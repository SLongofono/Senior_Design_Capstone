----------------------------------------------------------------------------------
-- Engineer: Longofono
-- 
-- Create Date: 11/13/2017 11:22:26 AM
-- Module Name: tb_decoder - Behavioral
-- Description: Test bench for decoder
-- 
-- Additional Comments:
-- 
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library config;
use work.config.all;

entity tb_decoder is
--  Port ( );
end tb_decoder;

architecture Behavioral of tb_decoder is

-- Components
component decode is
    Port(
        instr   : in std_logic_vector(63 downto 0);
        inst_t  : out instr_t;
        funct3  : out funct3_t;
        funct6  : out funct6_t;
        funct7  : out funct7_t;
        imm12   : out std_logic_vector(11 downto 0); -- I, B, and S Immediates
        imm20   : out std_logic_vector(20 downto 0); -- U and J Immediates
        opcode  : out opcode_t;
        rs1     : out reg_t;
        rs2     : out reg_t;
        rs3     : out reg_t;
        rd      : out reg_t;
        shamt   : out std_logic_vector(4 downto 0);
        csr     : out std_logic_vector(31 downto 20)
    );
end component;

-- Types for input
type test_input is array (0 to 157) of std_logic_vector(31 downto 0);

-- Signals
signal clk: std_logic := '0';
signal rst: std_logic := '1';
signal bin: std_logic_vector(31 downto 0) := (others => '0');
signal instr: instr_t;
signal s_funct3  : funct3_t;
signal s_funct6  : funct6_t;
signal s_funct7  : funct7_t;
signal s_imm12   : std_logic_vector(11 downto 0);
signal s_imm20   : std_logic_vector(20 downto 0);
signal s_opcode  : opcode_t;
signal s_rs1     : reg_t;
signal s_rs2     : reg_t;
signal s_rs3     : reg_t;
signal s_rd      : reg_t;
signal s_shamt   : std_logic_vector(4 downto 0);
signal s_csr     : std_logic_vector(31 downto 20)
signal inputs   : test_input :=
    (
    "00000000000000000000000000110111",
    "00000000000000000000000000010111",
    "00000000000000000000000001101111",
    "00000000000000000000000001100111",
    "00000000000000000000000001100011",
    "00000000000000000001000001100011",
    "00000000000000000100000001100011",
    "00000000000000000101000001100011",
    "00000000000000000110000001100011",
    "00000000000000000111000001100011",
    "00000000000000000000000000000011",
    "00000000000000000001000000000011",
    "00000000000000000010000000000011",
    "00000000000000000100000000000011",
    "00000000000000000101000000000011",
    "00000000000000000000000000100011",
    "00000000000000000001000000100011",
    "00000000000000000010000000100011",
    "00000000000000000000000000010011",
    "00000000000000000010000000010011",
    "00000000000000000011000000010011",
    "00000000000000000100000000010011",
    "00000000000000000110000000010011",
    "00000000000000000111000000010011",
    "00000000000000000001000000010011",
    "00000000000000000101000000010011",
    "01000000000000000101000000010011",
    "00000000000000000000000000110011",
    "01000000000000000000000000110011",
    "00000000000000000001000000110011",
    "00000000000000000010000000110011",
    "00000000000000000011000000110011",
    "00000000000000000100000000110011",
    "00000000000000000101000000110011",
    "01000000000000000101000000110011",
    "00000000000000000110000000110011",
    "00000000000000000111000000110011",
    "00000000000000000000000000001111",
    "00000000000000000001000000001111",
    "00000000000000000000000001110011",
    "00000000000100000000000001110011",
    "00000000000000000001000001110011",
    "00000000000000000010000001110011",
    "00000000000000000011000001110011",
    "00000000000000000101000001110011",
    "00000000000000000110000001110011",
    "00000000000000000111000001110011",
    "00000000000000000110000000000011",
    "00000000000000000011000000000011",
    "00000000000000000011000000100011",
    "00000000000000000001000000010011",
    "00000000000000000101000000010011",
    "01000000000000000101000000010011",
    "00000000000000000000000000011011",
    "00000000000000000001000000011011",
    "00000000000000000101000000011011",
    "01000000000000000101000000011011",
    "00000000000000000000000000111011",
    "01000000000000000000000000111011",
    "00000000000000000001000000111011",
    "00000000000000000101000000111011",
    "01000000000000000101000000111011",
    "00000010000000000000000000110011",
    "00000010000000000001000000110011",
    "00000010000000000010000000110011",
    "00000010000000000011000000110011",
    "00000010000000000100000000110011",
    "00000010000000000101000000110011",
    "00000010000000000110000000110011",
    "00000010000000000111000000110011",
    "00000010000000000000000000111011",
    "00000010000000000100000000111011",
    "00000010000000000101000000111011",
    "00000010000000000110000000111011",
    "00000010000000000111000000111011",
    "00010000000000000010000000101111",
    "00011000000000000010000000101111",
    "00001000000000000010000000101111",
    "00000000000000000010000000101111",
    "00100000000000000010000000101111",
    "01100000000000000010000000101111",
    "01000000000000000010000000101111",
    "10000000000000000010000000101111",
    "10100000000000000010000000101111",
    "11000000000000000010000000101111",
    "11100000000000000010000000101111",
    "00010000000000000011000000101111",
    "00011000000000000011000000101111",
    "00001000000000000011000000101111",
    "00000000000000000011000000101111",
    "00100000000000000011000000101111",
    "01100000000000000011000000101111",
    "01000000000000000011000000101111",
    "10000000000000000011000000101111",
    "10100000000000000011000000101111",
    "11000000000000000011000000101111",
    "11100000000000000011000000101111",
    "00000000000000000010000000000111",
    "00000000000000000010000000100111",
    "00000000000000000000000001000011",
    "00000000000000000000000001000111",
    "00000000000000000000000001001011",
    "00000000000000000000000001001111",
    "00000000000000000000000001010011",
    "00001000000000000000000001010011",
    "00010000000000000000000001010011",
    "00011000000000000000000001010011",
    "01011000000000000000000001010011",
    "00100000000000000000000001010011",
    "00100000000000000001000001010011",
    "00100000000000000010000001010011",
    "00101000000000000000000001010011",
    "00101000000000000001000001010011",
    "11000000000000000000000001010011",
    "11000000000100000000000001010011",
    "11100000000000000000000001010011",
    "10100000000000000010000001010011",
    "10100000000000000001000001010011",
    "10100000000000000000000001010011",
    "11100000000000000001000001010011",
    "11010000000000000000000001010011",
    "11010000000100000000000001010011",
    "11110000000000000000000001010011",
    "11000000001000000000000001010011",
    "11000000001100000000000001010011",
    "11010000001000000000000001010011",
    "11010000001100000000000001010011",
    "00000000000000000011000000000111",
    "00000000000000000011000000100111",
    "00000010000000000000000001000011",
    "00000010000000000000000001000111",
    "00000010000000000000000001001011",
    "00000010000000000000000001001111",
    "00000010000000000000000001010011",
    "00001010000000000000000001010011",
    "00010010000000000000000001010011",
    "00011010000000000000000001010011",
    "01011010000000000000000001010011",
    "00100010000000000000000001010011",
    "00100010000000000001000001010011",
    "00100010000000000010000001010011",
    "00101010000000000000000001010011",
    "00101010000000000001000001010011",
    "01000000000100000000000001010011",
    "01000010000000000000000001010011",
    "10100010000000000010000001010011",
    "10100010000000000001000001010011",
    "10100010000000000000000001010011",
    "11100010000000000001000001010011",
    "11000010000000000000000001010011",
    "11000010000100000000000001010011",
    "11010010000000000000000001010011",
    "11010010000100000000000001010011",
    "11000010001000000000000001010011",
    "11000010001100000000000001010011",
    "11100010000000000000000001010011",
    "11010010001000000000000001010011",
    "11010010001100000000000001010011",
    "11110010000000000000000001010011"
    );

begin

-- Declare components
dcode: decoder
    port map(
        instr => bin,
        inst_t => instr,
        funct3 => s_funct3,
        funct6 => s_funct6,
        funct7 => s_funct7,
        imm12 => s_imm12,
        imm20 => s_imm20,
        opcode => s_opcode,
        rs1 => s_rs1,
        rs2 => s_rs2,
        rs3 => s_rs3,
        rd => s_rd,
        shamt => s_shamt,
        csr => s_csr
    );

-- Clock generation
tiktok: process
begin
    wait for t_per/2;
    clk <= '0';
    wait for t_per/2;
    clk <= '1';
end process; -- end tiktok

main: process(clk)
begin
    wait for t_per;
    rst <= '0';
    
    for I in 0 to 157 loop
        bin <= inputs(I);
        wait for t_per;
    end loop;
    
    wait;
end process; --end main

end Behavioral;
