(0 + 0) => x"37", (0 + 1) => x"11", (0 + 2) => x"00", (0 + 3) => x"00", (0 + 4) => x"1b", (0 + 5) => x"01", (0 + 6) => x"71", (0 + 7) => x"80", (0 + 8) => x"13", (0 + 9) => x"11", (0 + 10) => x"41", (0 + 11) => x"01", (0 + 12) => x"6f", (0 + 13) => x"00", (0 + 14) => x"40", (0 + 15) => x"00", (0 + 16) => x"93", (0 + 17) => x"07", (0 + 18) => x"30", (0 + 19) => x"01", (0 + 20) => x"93", (0 + 21) => x"97", (0 + 22) => x"b7", (0 + 23) => x"01", (0 + 24) => x"13", (0 + 25) => x"07", (0 + 26) => x"10", (0 + 27) => x"00", (0 + 28) => x"23", (0 + 29) => x"90", (0 + 30) => x"e7", (0 + 31) => x"00", (0 + 32) => x"b7", (0 + 33) => x"17", (0 + 34) => x"80", (0 + 35) => x"09", (0 + 36) => x"97", (0 + 37) => x"06", (0 + 38) => x"00", (0 + 39) => x"00", (0 + 40) => x"93", (0 + 41) => x"86", (0 + 42) => x"46", (0 + 43) => x"09", (0 + 44) => x"13", (0 + 45) => x"07", (0 + 46) => x"10", (0 + 47) => x"02", (0 + 48) => x"93", (0 + 49) => x"97", (0 + 50) => x"47", (0 + 51) => x"00", (0 + 52) => x"93", (0 + 53) => x"05", (0 + 54) => x"10", (0 + 55) => x"00", (0 + 56) => x"03", (0 + 57) => x"c6", (0 + 58) => x"47", (0 + 59) => x"00", (0 + 60) => x"13", (0 + 61) => x"76", (0 + 62) => x"f6", (0 + 63) => x"0f", (0 + 64) => x"e3", (0 + 65) => x"0c", (0 + 66) => x"06", (0 + 67) => x"fe", (0 + 68) => x"a3", (0 + 69) => x"81", (0 + 70) => x"e7", (0 + 71) => x"00", (0 + 72) => x"a3", (0 + 73) => x"82", (0 + 74) => x"b7", (0 + 75) => x"00", (0 + 76) => x"93", (0 + 77) => x"86", (0 + 78) => x"16", (0 + 79) => x"00", (0 + 80) => x"03", (0 + 81) => x"c7", (0 + 82) => x"06", (0 + 83) => x"00", (0 + 84) => x"e3", (0 + 85) => x"12", (0 + 86) => x"07", (0 + 87) => x"fe", (0 + 88) => x"37", (0 + 89) => x"17", (0 + 90) => x"80", (0 + 91) => x"09", (0 + 92) => x"13", (0 + 93) => x"05", (0 + 94) => x"30", (0 + 95) => x"01", (0 + 96) => x"93", (0 + 97) => x"06", (0 + 98) => x"10", (0 + 99) => x"00", (0 + 100) => x"13", (0 + 101) => x"17", (0 + 102) => x"47", (0 + 103) => x"00", (0 + 104) => x"93", (0 + 105) => x"05", (0 + 106) => x"10", (0 + 107) => x"00", (0 + 108) => x"13", (0 + 109) => x"15", (0 + 110) => x"b5", (0 + 111) => x"01", (0 + 112) => x"83", (0 + 113) => x"47", (0 + 114) => x"17", (0 + 115) => x"00", (0 + 116) => x"93", (0 + 117) => x"f7", (0 + 118) => x"f7", (0 + 119) => x"0f", (0 + 120) => x"e3", (0 + 121) => x"8c", (0 + 122) => x"07", (0 + 123) => x"fe", (0 + 124) => x"03", (0 + 125) => x"46", (0 + 126) => x"07", (0 + 127) => x"00", (0 + 128) => x"9b", (0 + 129) => x"86", (0 + 130) => x"16", (0 + 131) => x"00", (0 + 132) => x"93", (0 + 133) => x"96", (0 + 134) => x"06", (0 + 135) => x"03", (0 + 136) => x"23", (0 + 137) => x"01", (0 + 138) => x"b7", (0 + 139) => x"00", (0 + 140) => x"93", (0 + 141) => x"d6", (0 + 142) => x"06", (0 + 143) => x"03", (0 + 144) => x"13", (0 + 145) => x"76", (0 + 146) => x"f6", (0 + 147) => x"0f", (0 + 148) => x"23", (0 + 149) => x"10", (0 + 150) => x"d5", (0 + 151) => x"00", (0 + 152) => x"83", (0 + 153) => x"47", (0 + 154) => x"47", (0 + 155) => x"00", (0 + 156) => x"93", (0 + 157) => x"f7", (0 + 158) => x"f7", (0 + 159) => x"0f", (0 + 160) => x"e3", (0 + 161) => x"8c", (0 + 162) => x"07", (0 + 163) => x"fe", (0 + 164) => x"a3", (0 + 165) => x"01", (0 + 166) => x"c7", (0 + 167) => x"00", (0 + 168) => x"a3", (0 + 169) => x"02", (0 + 170) => x"b7", (0 + 171) => x"00", (0 + 172) => x"6f", (0 + 173) => x"f0", (0 + 174) => x"5f", (0 + 175) => x"fc", (0 + 176) => x"00", (0 + 177) => x"00", (0 + 178) => x"00", (0 + 179) => x"00", (0 + 180) => x"00", (0 + 181) => x"00", (0 + 182) => x"00", (0 + 183) => x"00", (0 + 184) => x"21", (0 + 185) => x"21", (0 + 186) => x"21", (0 + 187) => x"45", (0 + 188) => x"43", (0 + 189) => x"48", (0 + 190) => x"4f", (0 + 191) => x"20", (0 + 192) => x"53", (0 + 193) => x"45", (0 + 194) => x"52", (0 + 195) => x"56", (0 + 196) => x"45", (0 + 197) => x"52", (0 + 198) => x"21", (0 + 199) => x"21", (0 + 200) => x"21", (0 + 201) => x"0a", (0 + 202) => x"00", (0 + 203) => x"00", (0 + 204) => x"00", (0 + 205) => x"00", (0 + 206) => x"00", (0 + 207) => x"00", (0 + 208) => x"00", (0 + 209) => x"00", (0 + 210) => x"00", (0 + 211) => x"00", (0 + 212) => x"00", (0 + 213) => x"00", (0 + 214) => x"00", (0 + 215) => x"00", (0 + 216) => x"00", (0 + 217) => x"00", (0 + 218) => x"00", (0 + 219) => x"00", (0 + 220) => x"00", (0 + 221) => x"00", (0 + 222) => x"00", (0 + 223) => x"00", (0 + 224) => x"00", (0 + 225) => x"00", (0 + 226) => x"00", (0 + 227) => x"00", (0 + 228) => x"00", (0 + 229) => x"00", (0 + 230) => x"00", (0 + 231) => x"00", (0 + 232) => x"00", (0 + 233) => x"00", (0 + 234) => x"00", (0 + 235) => x"00", (0 + 236) => x"00", (0 + 237) => x"00", (0 + 238) => x"00", (0 + 239) => x"00", (0 + 240) => x"00", (0 + 241) => x"00", (0 + 242) => x"00", (0 + 243) => x"00", (0 + 244) => x"00", (0 + 245) => x"00", (0 + 246) => x"00", (0 + 247) => x"00", (0 + 248) => x"00", (0 + 249) => x"00", (0 + 250) => x"00", (0 + 251) => x"00", (0 + 252) => x"00", (0 + 253) => x"00", (0 + 254) => x"00", (0 + 255) => x"00", (0 + 256) => x"00", (0 + 257) => x"00", (0 + 258) => x"00", (0 + 259) => x"00", (0 + 260) => x"00", (0 + 261) => x"00", (0 + 262) => x"00", (0 + 263) => x"00", (0 + 264) => x"00", (0 + 265) => x"00", (0 + 266) => x"00", (0 + 267) => x"00", (0 + 268) => x"00", (0 + 269) => x"00", (0 + 270) => x"00", (0 + 271) => x"00", (0 + 272) => x"00", (0 + 273) => x"00", (0 + 274) => x"00", (0 + 275) => x"00", (0 + 276) => x"00", (0 + 277) => x"00", (0 + 278) => x"00", (0 + 279) => x"00", (0 + 280) => x"00", (0 + 281) => x"00", (0 + 282) => x"00", (0 + 283) => x"00", (0 + 284) => x"00", (0 + 285) => x"00", (0 + 286) => x"00", (0 + 287) => x"00", (0 + 288) => x"00", (0 + 289) => x"00", (0 + 290) => x"00", (0 + 291) => x"00", (0 + 292) => x"00", (0 + 293) => x"00", (0 + 294) => x"00", (0 + 295) => x"00", (0 + 296) => x"00", (0 + 297) => x"00", (0 + 298) => x"00", (0 + 299) => x"00", (0 + 300) => x"00", (0 + 301) => x"00", (0 + 302) => x"00", (0 + 303) => x"00", (0 + 304) => x"00", (0 + 305) => x"00", (0 + 306) => x"00", (0 + 307) => x"00", (0 + 308) => x"00", (0 + 309) => x"00", (0 + 310) => x"00", (0 + 311) => x"00", (0 + 312) => x"00", (0 + 313) => x"00", (0 + 314) => x"00", (0 + 315) => x"00", (0 + 316) => x"00", (0 + 317) => x"00", (0 + 318) => x"00", (0 + 319) => x"00", (0 + 320) => x"00", (0 + 321) => x"00", (0 + 322) => x"00", (0 + 323) => x"00", (0 + 324) => x"00", (0 + 325) => x"00", (0 + 326) => x"00", (0 + 327) => x"00", (0 + 328) => x"00", (0 + 329) => x"00", (0 + 330) => x"00", (0 + 331) => x"00", (0 + 332) => x"00", (0 + 333) => x"00", (0 + 334) => x"00", (0 + 335) => x"00", (0 + 336) => x"00", (0 + 337) => x"00", (0 + 338) => x"00", (0 + 339) => x"00", (0 + 340) => x"00", (0 + 341) => x"00", (0 + 342) => x"00", (0 + 343) => x"00", (0 + 344) => x"00", (0 + 345) => x"00", (0 + 346) => x"00", (0 + 347) => x"00", (0 + 348) => x"00", (0 + 349) => x"00", (0 + 350) => x"00", (0 + 351) => x"00", (0 + 352) => x"00", (0 + 353) => x"00", (0 + 354) => x"00", (0 + 355) => x"00", (0 + 356) => x"00", (0 + 357) => x"00", (0 + 358) => x"00", (0 + 359) => x"00", (0 + 360) => x"00", (0 + 361) => x"00", (0 + 362) => x"00", (0 + 363) => x"00", (0 + 364) => x"00", (0 + 365) => x"00", (0 + 366) => x"00", (0 + 367) => x"00", (0 + 368) => x"00", (0 + 369) => x"00", (0 + 370) => x"00", (0 + 371) => x"00", (0 + 372) => x"00", (0 + 373) => x"00", (0 + 374) => x"00", (0 + 375) => x"00", (0 + 376) => x"00", (0 + 377) => x"00", (0 + 378) => x"00", (0 + 379) => x"00", (0 + 380) => x"00", (0 + 381) => x"00", (0 + 382) => x"00", (0 + 383) => x"00", (0 + 384) => x"00", (0 + 385) => x"00", (0 + 386) => x"00", (0 + 387) => x"00", (0 + 388) => x"00", (0 + 389) => x"00", (0 + 390) => x"00", (0 + 391) => x"00", (0 + 392) => x"00", (0 + 393) => x"00", (0 + 394) => x"00", (0 + 395) => x"00", (0 + 396) => x"00", (0 + 397) => x"00", (0 + 398) => x"00", (0 + 399) => x"00", (0 + 400) => x"00", (0 + 401) => x"00", (0 + 402) => x"00", (0 + 403) => x"00", (0 + 404) => x"00", (0 + 405) => x"00", (0 + 406) => x"00", (0 + 407) => x"00", (0 + 408) => x"00", (0 + 409) => x"00", (0 + 410) => x"00", (0 + 411) => x"00", (0 + 412) => x"00", (0 + 413) => x"00", (0 + 414) => x"00", (0 + 415) => x"00", (0 + 416) => x"00", (0 + 417) => x"00", (0 + 418) => x"00", (0 + 419) => x"00", (0 + 420) => x"00", (0 + 421) => x"00", (0 + 422) => x"00", (0 + 423) => x"00", (0 + 424) => x"00", (0 + 425) => x"00", (0 + 426) => x"00", (0 + 427) => x"00", (0 + 428) => x"00", (0 + 429) => x"00", (0 + 430) => x"00", (0 + 431) => x"00", (0 + 432) => x"00", (0 + 433) => x"00", (0 + 434) => x"00", (0 + 435) => x"00", (0 + 436) => x"00", (0 + 437) => x"00", (0 + 438) => x"00", (0 + 439) => x"00", (0 + 440) => x"00", (0 + 441) => x"00", (0 + 442) => x"00", (0 + 443) => x"00", (0 + 444) => x"00", (0 + 445) => x"00", (0 + 446) => x"00", (0 + 447) => x"00", (0 + 448) => x"00", (0 + 449) => x"00", (0 + 450) => x"00", (0 + 451) => x"00", (0 + 452) => x"00", (0 + 453) => x"00", (0 + 454) => x"00", (0 + 455) => x"00", (0 + 456) => x"00", (0 + 457) => x"00", (0 + 458) => x"00", (0 + 459) => x"00", (0 + 460) => x"00", (0 + 461) => x"00", (0 + 462) => x"00", (0 + 463) => x"00", (0 + 464) => x"00", (0 + 465) => x"00", (0 + 466) => x"00", (0 + 467) => x"00", (0 + 468) => x"00", (0 + 469) => x"00", (0 + 470) => x"00", (0 + 471) => x"00", (0 + 472) => x"00", (0 + 473) => x"00", (0 + 474) => x"00", (0 + 475) => x"00", (0 + 476) => x"00", (0 + 477) => x"00", (0 + 478) => x"00", (0 + 479) => x"00", (0 + 480) => x"00", (0 + 481) => x"00", (0 + 482) => x"00", (0 + 483) => x"00", (0 + 484) => x"00", (0 + 485) => x"00", (0 + 486) => x"00", (0 + 487) => x"00", (0 + 488) => x"00", (0 + 489) => x"00", (0 + 490) => x"00", (0 + 491) => x"00", (0 + 492) => x"00", (0 + 493) => x"00", (0 + 494) => x"00", (0 + 495) => x"00", (0 + 496) => x"00", (0 + 497) => x"00", (0 + 498) => x"00", (0 + 499) => x"00", (0 + 500) => x"00", (0 + 501) => x"00", (0 + 502) => x"00", (0 + 503) => x"00", (0 + 504) => x"00", (0 + 505) => x"00", (0 + 506) => x"00", (0 + 507) => x"00", (0 + 508) => x"00", (0 + 509) => x"00", (0 + 510) => x"00", (0 + 511) => x"00", (0 + 512) => x"00", (0 + 513) => x"00", (0 + 514) => x"00", (0 + 515) => x"00", (0 + 516) => x"00", (0 + 517) => x"00", (0 + 518) => x"00", (0 + 519) => x"00", (0 + 520) => x"00", (0 + 521) => x"00", (0 + 522) => x"00", (0 + 523) => x"00", (0 + 524) => x"00", (0 + 525) => x"00", (0 + 526) => x"00", (0 + 527) => x"00", (0 + 528) => x"00", (0 + 529) => x"00", (0 + 530) => x"00", (0 + 531) => x"00", (0 + 532) => x"00", (0 + 533) => x"00", (0 + 534) => x"00", (0 + 535) => x"00", (0 + 536) => x"00", (0 + 537) => x"00", (0 + 538) => x"00", (0 + 539) => x"00", (0 + 540) => x"00", (0 + 541) => x"00", (0 + 542) => x"00", (0 + 543) => x"00", (0 + 544) => x"00", (0 + 545) => x"00", (0 + 546) => x"00", (0 + 547) => x"00", (0 + 548) => x"00", (0 + 549) => x"00", (0 + 550) => x"00", (0 + 551) => x"00", (0 + 552) => x"00", (0 + 553) => x"00", (0 + 554) => x"00", (0 + 555) => x"00", (0 + 556) => x"00", (0 + 557) => x"00", (0 + 558) => x"00", (0 + 559) => x"00", (0 + 560) => x"00", (0 + 561) => x"00", (0 + 562) => x"00", (0 + 563) => x"00", (0 + 564) => x"00", (0 + 565) => x"00", (0 + 566) => x"00", (0 + 567) => x"00", (0 + 568) => x"00", (0 + 569) => x"00", (0 + 570) => x"00", (0 + 571) => x"00", (0 + 572) => x"00", (0 + 573) => x"00", (0 + 574) => x"00", (0 + 575) => x"00", (0 + 576) => x"00", (0 + 577) => x"00", (0 + 578) => x"00", (0 + 579) => x"00", (0 + 580) => x"00", (0 + 581) => x"00", (0 + 582) => x"00", (0 + 583) => x"00", (0 + 584) => x"00", (0 + 585) => x"00", (0 + 586) => x"00", (0 + 587) => x"00", (0 + 588) => x"00", (0 + 589) => x"00", (0 + 590) => x"00", (0 + 591) => x"00", (0 + 592) => x"00", (0 + 593) => x"00", (0 + 594) => x"00", (0 + 595) => x"00", (0 + 596) => x"00", (0 + 597) => x"00", (0 + 598) => x"00", (0 + 599) => x"00", (0 + 600) => x"00", (0 + 601) => x"00", (0 + 602) => x"00", (0 + 603) => x"00", (0 + 604) => x"00", (0 + 605) => x"00", (0 + 606) => x"00", (0 + 607) => x"00", (0 + 608) => x"00", (0 + 609) => x"00", (0 + 610) => x"00", (0 + 611) => x"00", (0 + 612) => x"00", (0 + 613) => x"00", (0 + 614) => x"00", (0 + 615) => x"00", (0 + 616) => x"00", (0 + 617) => x"00", (0 + 618) => x"00", (0 + 619) => x"00", (0 + 620) => x"00", (0 + 621) => x"00", (0 + 622) => x"00", (0 + 623) => x"00", (0 + 624) => x"00", (0 + 625) => x"00", (0 + 626) => x"00", (0 + 627) => x"00", (0 + 628) => x"00", (0 + 629) => x"00", (0 + 630) => x"00", (0 + 631) => x"00", (0 + 632) => x"00", (0 + 633) => x"00", (0 + 634) => x"00", (0 + 635) => x"00", (0 + 636) => x"00", (0 + 637) => x"00", (0 + 638) => x"00", (0 + 639) => x"00", (0 + 640) => x"00", (0 + 641) => x"00", (0 + 642) => x"00", (0 + 643) => x"00", (0 + 644) => x"00", (0 + 645) => x"00", (0 + 646) => x"00", (0 + 647) => x"00", (0 + 648) => x"00", (0 + 649) => x"00", (0 + 650) => x"00", (0 + 651) => x"00", (0 + 652) => x"00", (0 + 653) => x"00", (0 + 654) => x"00", (0 + 655) => x"00", (0 + 656) => x"00", (0 + 657) => x"00", (0 + 658) => x"00", (0 + 659) => x"00", (0 + 660) => x"00", (0 + 661) => x"00", (0 + 662) => x"00", (0 + 663) => x"00", (0 + 664) => x"00", (0 + 665) => x"00", (0 + 666) => x"00", (0 + 667) => x"00", (0 + 668) => x"00", (0 + 669) => x"00", (0 + 670) => x"00", (0 + 671) => x"00", (0 + 672) => x"00", (0 + 673) => x"00", (0 + 674) => x"00", (0 + 675) => x"00", (0 + 676) => x"00", (0 + 677) => x"00", (0 + 678) => x"00", (0 + 679) => x"00", (0 + 680) => x"00", (0 + 681) => x"00", (0 + 682) => x"00", (0 + 683) => x"00", (0 + 684) => x"00", (0 + 685) => x"00", (0 + 686) => x"00", (0 + 687) => x"00", (0 + 688) => x"00", (0 + 689) => x"00", (0 + 690) => x"00", (0 + 691) => x"00", (0 + 692) => x"00", (0 + 693) => x"00", (0 + 694) => x"00", (0 + 695) => x"00", (0 + 696) => x"00", (0 + 697) => x"00", (0 + 698) => x"00", (0 + 699) => x"00", (0 + 700) => x"00", (0 + 701) => x"00", (0 + 702) => x"00", (0 + 703) => x"00", (0 + 704) => x"00", (0 + 705) => x"00", (0 + 706) => x"00", (0 + 707) => x"00", (0 + 708) => x"00", (0 + 709) => x"00", (0 + 710) => x"00", (0 + 711) => x"00", (0 + 712) => x"00", (0 + 713) => x"00", (0 + 714) => x"00", (0 + 715) => x"00", (0 + 716) => x"00", (0 + 717) => x"00", (0 + 718) => x"00", (0 + 719) => x"00", (0 + 720) => x"00", (0 + 721) => x"00", (0 + 722) => x"00", (0 + 723) => x"00", (0 + 724) => x"00", (0 + 725) => x"00", (0 + 726) => x"00", (0 + 727) => x"00", (0 + 728) => x"00", (0 + 729) => x"00", (0 + 730) => x"00", (0 + 731) => x"00", (0 + 732) => x"00", (0 + 733) => x"00", (0 + 734) => x"00", (0 + 735) => x"00", (0 + 736) => x"00", (0 + 737) => x"00", (0 + 738) => x"00", (0 + 739) => x"00", (0 + 740) => x"00", (0 + 741) => x"00", (0 + 742) => x"00", (0 + 743) => x"00", (0 + 744) => x"00", (0 + 745) => x"00", (0 + 746) => x"00", (0 + 747) => x"00", (0 + 748) => x"00", (0 + 749) => x"00", (0 + 750) => x"00", (0 + 751) => x"00", (0 + 752) => x"00", (0 + 753) => x"00", (0 + 754) => x"00", (0 + 755) => x"00", (0 + 756) => x"00", (0 + 757) => x"00", (0 + 758) => x"00", (0 + 759) => x"00", (0 + 760) => x"00", (0 + 761) => x"00", (0 + 762) => x"00", (0 + 763) => x"00", (0 + 764) => x"00", (0 + 765) => x"00", (0 + 766) => x"00", (0 + 767) => x"00", (0 + 768) => x"00", (0 + 769) => x"00", (0 + 770) => x"00", (0 + 771) => x"00", (0 + 772) => x"00", (0 + 773) => x"00", (0 + 774) => x"00", (0 + 775) => x"00", (0 + 776) => x"00", (0 + 777) => x"00", (0 + 778) => x"00", (0 + 779) => x"00", (0 + 780) => x"00", (0 + 781) => x"00", (0 + 782) => x"00", (0 + 783) => x"00", (0 + 784) => x"00", (0 + 785) => x"00", (0 + 786) => x"00", (0 + 787) => x"00", (0 + 788) => x"00", (0 + 789) => x"00", (0 + 790) => x"00", (0 + 791) => x"00", (0 + 792) => x"00", (0 + 793) => x"00", (0 + 794) => x"00", (0 + 795) => x"00", (0 + 796) => x"00", (0 + 797) => x"00", (0 + 798) => x"00", (0 + 799) => x"00", (0 + 800) => x"00", (0 + 801) => x"00", (0 + 802) => x"00", (0 + 803) => x"00", (0 + 804) => x"00", (0 + 805) => x"00", (0 + 806) => x"00", (0 + 807) => x"00", (0 + 808) => x"00", (0 + 809) => x"00", (0 + 810) => x"00", (0 + 811) => x"00", (0 + 812) => x"00", (0 + 813) => x"00", (0 + 814) => x"00", (0 + 815) => x"00", (0 + 816) => x"00", (0 + 817) => x"00", (0 + 818) => x"00", (0 + 819) => x"00", (0 + 820) => x"00", (0 + 821) => x"00", (0 + 822) => x"00", (0 + 823) => x"00", (0 + 824) => x"00", (0 + 825) => x"00", (0 + 826) => x"00", (0 + 827) => x"00", (0 + 828) => x"00", (0 + 829) => x"00", (0 + 830) => x"00", (0 + 831) => x"00", (0 + 832) => x"00", (0 + 833) => x"00", (0 + 834) => x"00", (0 + 835) => x"00", (0 + 836) => x"00", (0 + 837) => x"00", (0 + 838) => x"00", (0 + 839) => x"00", (0 + 840) => x"00", (0 + 841) => x"00", (0 + 842) => x"00", (0 + 843) => x"00", (0 + 844) => x"00", (0 + 845) => x"00", (0 + 846) => x"00", (0 + 847) => x"00", (0 + 848) => x"00", (0 + 849) => x"00", (0 + 850) => x"00", (0 + 851) => x"00", (0 + 852) => x"00", (0 + 853) => x"00", (0 + 854) => x"00", (0 + 855) => x"00", (0 + 856) => x"00", (0 + 857) => x"00", (0 + 858) => x"00", (0 + 859) => x"00", (0 + 860) => x"00", (0 + 861) => x"00", (0 + 862) => x"00", (0 + 863) => x"00", (0 + 864) => x"00", (0 + 865) => x"00", (0 + 866) => x"00", (0 + 867) => x"00", (0 + 868) => x"00", (0 + 869) => x"00", (0 + 870) => x"00", (0 + 871) => x"00", (0 + 872) => x"00", (0 + 873) => x"00", (0 + 874) => x"00", (0 + 875) => x"00", (0 + 876) => x"00", (0 + 877) => x"00", (0 + 878) => x"00", (0 + 879) => x"00", (0 + 880) => x"00", (0 + 881) => x"00", (0 + 882) => x"00", (0 + 883) => x"00", (0 + 884) => x"00", (0 + 885) => x"00", (0 + 886) => x"00", (0 + 887) => x"00", (0 + 888) => x"00", (0 + 889) => x"00", (0 + 890) => x"00", (0 + 891) => x"00", (0 + 892) => x"00", (0 + 893) => x"00", (0 + 894) => x"00", (0 + 895) => x"00", (0 + 896) => x"00", (0 + 897) => x"00", (0 + 898) => x"00", (0 + 899) => x"00", (0 + 900) => x"00", (0 + 901) => x"00", (0 + 902) => x"00", (0 + 903) => x"00", (0 + 904) => x"00", (0 + 905) => x"00", (0 + 906) => x"00", (0 + 907) => x"00", (0 + 908) => x"00", (0 + 909) => x"00", (0 + 910) => x"00", (0 + 911) => x"00", (0 + 912) => x"00", (0 + 913) => x"00", (0 + 914) => x"00", (0 + 915) => x"00", (0 + 916) => x"00", (0 + 917) => x"00", (0 + 918) => x"00", (0 + 919) => x"00", (0 + 920) => x"00", (0 + 921) => x"00", (0 + 922) => x"00", (0 + 923) => x"00", (0 + 924) => x"00", (0 + 925) => x"00", (0 + 926) => x"00", (0 + 927) => x"00", (0 + 928) => x"00", (0 + 929) => x"00", (0 + 930) => x"00", (0 + 931) => x"00", (0 + 932) => x"00", (0 + 933) => x"00", (0 + 934) => x"00", (0 + 935) => x"00", (0 + 936) => x"00", (0 + 937) => x"00", (0 + 938) => x"00", (0 + 939) => x"00", (0 + 940) => x"00", (0 + 941) => x"00", (0 + 942) => x"00", (0 + 943) => x"00", (0 + 944) => x"00", (0 + 945) => x"00", (0 + 946) => x"00", (0 + 947) => x"00", (0 + 948) => x"00", (0 + 949) => x"00", (0 + 950) => x"00", (0 + 951) => x"00", (0 + 952) => x"00", (0 + 953) => x"00", (0 + 954) => x"00", (0 + 955) => x"00", (0 + 956) => x"00", (0 + 957) => x"00", (0 + 958) => x"00", (0 + 959) => x"00", (0 + 960) => x"00", (0 + 961) => x"00", (0 + 962) => x"00", (0 + 963) => x"00", (0 + 964) => x"00", (0 + 965) => x"00", (0 + 966) => x"00", (0 + 967) => x"00", (0 + 968) => x"00", (0 + 969) => x"00", (0 + 970) => x"00", (0 + 971) => x"00", (0 + 972) => x"00", (0 + 973) => x"00", (0 + 974) => x"00", (0 + 975) => x"00", (0 + 976) => x"00", (0 + 977) => x"00", (0 + 978) => x"00", (0 + 979) => x"00", (0 + 980) => x"00", (0 + 981) => x"00", (0 + 982) => x"00", (0 + 983) => x"00", (0 + 984) => x"00", (0 + 985) => x"00", (0 + 986) => x"00", (0 + 987) => x"00", (0 + 988) => x"00", (0 + 989) => x"00", (0 + 990) => x"00", (0 + 991) => x"00", (0 + 992) => x"00", (0 + 993) => x"00", (0 + 994) => x"00", (0 + 995) => x"00", (0 + 996) => x"00", (0 + 997) => x"00", (0 + 998) => x"00", (0 + 999) => x"00", (0 + 1000) => x"00", (0 + 1001) => x"00", (0 + 1002) => x"00", (0 + 1003) => x"00", (0 + 1004) => x"00", (0 + 1005) => x"00", (0 + 1006) => x"00", (0 + 1007) => x"00", (0 + 1008) => x"00", (0 + 1009) => x"00", (0 + 1010) => x"00", (0 + 1011) => x"00", (0 + 1012) => x"00", (0 + 1013) => x"00", (0 + 1014) => x"00", (0 + 1015) => x"00", (0 + 1016) => x"00", (0 + 1017) => x"00", (0 + 1018) => x"00", (0 + 1019) => x"00", (0 + 1020) => x"00", (0 + 1021) => x"00", (0 + 1022) => x"00", (0 + 1023) => x"00", (0 + 1024) => x"00", (0 + 1025) => x"00", (0 + 1026) => x"00", (0 + 1027) => x"00", (0 + 1028) => x"00", (0 + 1029) => x"00", (0 + 1030) => x"00", (0 + 1031) => x"00", (0 + 1032) => x"00", (0 + 1033) => x"00", (0 + 1034) => x"00", (0 + 1035) => x"00", (0 + 1036) => x"00", (0 + 1037) => x"00", (0 + 1038) => x"00", (0 + 1039) => x"00", (0 + 1040) => x"00", (0 + 1041) => x"00", (0 + 1042) => x"00", (0 + 1043) => x"00", (0 + 1044) => x"00", (0 + 1045) => x"00", (0 + 1046) => x"00", (0 + 1047) => x"00", (0 + 1048) => x"00", (0 + 1049) => x"00", (0 + 1050) => x"00", (0 + 1051) => x"00", (0 + 1052) => x"00", (0 + 1053) => x"00", (0 + 1054) => x"00", (0 + 1055) => x"00", (0 + 1056) => x"00", (0 + 1057) => x"00", (0 + 1058) => x"00", (0 + 1059) => x"00", (0 + 1060) => x"00", (0 + 1061) => x"00", (0 + 1062) => x"00", (0 + 1063) => x"00", (0 + 1064) => x"00", (0 + 1065) => x"00", (0 + 1066) => x"00", (0 + 1067) => x"00", (0 + 1068) => x"00", (0 + 1069) => x"00", (0 + 1070) => x"00", (0 + 1071) => x"00", (0 + 1072) => x"00", (0 + 1073) => x"00", (0 + 1074) => x"00", (0 + 1075) => x"00", (0 + 1076) => x"00", (0 + 1077) => x"00", (0 + 1078) => x"00", (0 + 1079) => x"00", (0 + 1080) => x"00", (0 + 1081) => x"00", (0 + 1082) => x"00", (0 + 1083) => x"00", (0 + 1084) => x"00", (0 + 1085) => x"00", (0 + 1086) => x"00", (0 + 1087) => x"00", (0 + 1088) => x"00", (0 + 1089) => x"00", (0 + 1090) => x"00", (0 + 1091) => x"00", (0 + 1092) => x"00", (0 + 1093) => x"00", (0 + 1094) => x"00", (0 + 1095) => x"00", (0 + 1096) => x"00", (0 + 1097) => x"00", (0 + 1098) => x"00", (0 + 1099) => x"00", (0 + 1100) => x"00", (0 + 1101) => x"00", (0 + 1102) => x"00", (0 + 1103) => x"00", (0 + 1104) => x"00", (0 + 1105) => x"00", (0 + 1106) => x"00", (0 + 1107) => x"00", (0 + 1108) => x"00", (0 + 1109) => x"00", (0 + 1110) => x"00", (0 + 1111) => x"00", (0 + 1112) => x"00", (0 + 1113) => x"00", (0 + 1114) => x"00", (0 + 1115) => x"00", (0 + 1116) => x"00", (0 + 1117) => x"00", (0 + 1118) => x"00", (0 + 1119) => x"00", (0 + 1120) => x"00", (0 + 1121) => x"00", (0 + 1122) => x"00", (0 + 1123) => x"00", (0 + 1124) => x"00", (0 + 1125) => x"00", (0 + 1126) => x"00", (0 + 1127) => x"00", (0 + 1128) => x"00", (0 + 1129) => x"00", (0 + 1130) => x"00", (0 + 1131) => x"00", (0 + 1132) => x"00", (0 + 1133) => x"00", (0 + 1134) => x"00", (0 + 1135) => x"00", (0 + 1136) => x"00", (0 + 1137) => x"00", (0 + 1138) => x"00", (0 + 1139) => x"00", (0 + 1140) => x"00", (0 + 1141) => x"00", (0 + 1142) => x"00", (0 + 1143) => x"00", (0 + 1144) => x"00", (0 + 1145) => x"00", (0 + 1146) => x"00", (0 + 1147) => x"00", (0 + 1148) => x"00", (0 + 1149) => x"00", (0 + 1150) => x"00", (0 + 1151) => x"00", (0 + 1152) => x"00", (0 + 1153) => x"00", (0 + 1154) => x"00", (0 + 1155) => x"00", (0 + 1156) => x"00", (0 + 1157) => x"00", (0 + 1158) => x"00", (0 + 1159) => x"00", (0 + 1160) => x"00", (0 + 1161) => x"00", (0 + 1162) => x"00", (0 + 1163) => x"00", (0 + 1164) => x"00", (0 + 1165) => x"00", (0 + 1166) => x"00", (0 + 1167) => x"00", (0 + 1168) => x"00", (0 + 1169) => x"00", (0 + 1170) => x"00", (0 + 1171) => x"00", (0 + 1172) => x"00", (0 + 1173) => x"00", (0 + 1174) => x"00", (0 + 1175) => x"00", (0 + 1176) => x"00", (0 + 1177) => x"00", (0 + 1178) => x"00", (0 + 1179) => x"00", (0 + 1180) => x"00", (0 + 1181) => x"00", (0 + 1182) => x"00", (0 + 1183) => x"00", (0 + 1184) => x"00", (0 + 1185) => x"00", (0 + 1186) => x"00", (0 + 1187) => x"00", (0 + 1188) => x"00", (0 + 1189) => x"00", (0 + 1190) => x"00", (0 + 1191) => x"00", (0 + 1192) => x"00", (0 + 1193) => x"00", (0 + 1194) => x"00", (0 + 1195) => x"00", (0 + 1196) => x"00", (0 + 1197) => x"00", (0 + 1198) => x"00", (0 + 1199) => x"00", (0 + 1200) => x"00", (0 + 1201) => x"00", (0 + 1202) => x"00", (0 + 1203) => x"00", (0 + 1204) => x"00", (0 + 1205) => x"00", (0 + 1206) => x"00", (0 + 1207) => x"00", (0 + 1208) => x"00", (0 + 1209) => x"00", (0 + 1210) => x"00", (0 + 1211) => x"00", (0 + 1212) => x"00", (0 + 1213) => x"00", (0 + 1214) => x"00", (0 + 1215) => x"00", (0 + 1216) => x"00", (0 + 1217) => x"00", (0 + 1218) => x"00", (0 + 1219) => x"00", (0 + 1220) => x"00", (0 + 1221) => x"00", (0 + 1222) => x"00", (0 + 1223) => x"00", (0 + 1224) => x"00", (0 + 1225) => x"00", (0 + 1226) => x"00", (0 + 1227) => x"00", (0 + 1228) => x"00", (0 + 1229) => x"00", (0 + 1230) => x"00", (0 + 1231) => x"00", (0 + 1232) => x"00", (0 + 1233) => x"00", (0 + 1234) => x"00", (0 + 1235) => x"00", (0 + 1236) => x"00", (0 + 1237) => x"00", (0 + 1238) => x"00", (0 + 1239) => x"00", (0 + 1240) => x"00", (0 + 1241) => x"00", (0 + 1242) => x"00", (0 + 1243) => x"00", (0 + 1244) => x"00", (0 + 1245) => x"00", (0 + 1246) => x"00", (0 + 1247) => x"00", (0 + 1248) => x"00", (0 + 1249) => x"00", (0 + 1250) => x"00", (0 + 1251) => x"00", (0 + 1252) => x"00", (0 + 1253) => x"00", (0 + 1254) => x"00", (0 + 1255) => x"00", (0 + 1256) => x"00", (0 + 1257) => x"00", (0 + 1258) => x"00", (0 + 1259) => x"00", (0 + 1260) => x"00", (0 + 1261) => x"00", (0 + 1262) => x"00", (0 + 1263) => x"00", (0 + 1264) => x"00", (0 + 1265) => x"00", (0 + 1266) => x"00", (0 + 1267) => x"00", (0 + 1268) => x"00", (0 + 1269) => x"00", (0 + 1270) => x"00", (0 + 1271) => x"00", (0 + 1272) => x"00", (0 + 1273) => x"00", (0 + 1274) => x"00", (0 + 1275) => x"00", (0 + 1276) => x"00", (0 + 1277) => x"00", (0 + 1278) => x"00", (0 + 1279) => x"00", (0 + 1280) => x"00", (0 + 1281) => x"00", (0 + 1282) => x"00", (0 + 1283) => x"00", (0 + 1284) => x"00", (0 + 1285) => x"00", (0 + 1286) => x"00", (0 + 1287) => x"00", (0 + 1288) => x"00", (0 + 1289) => x"00", (0 + 1290) => x"00", (0 + 1291) => x"00", (0 + 1292) => x"00", (0 + 1293) => x"00", (0 + 1294) => x"00", (0 + 1295) => x"00", (0 + 1296) => x"00", (0 + 1297) => x"00", (0 + 1298) => x"00", (0 + 1299) => x"00", (0 + 1300) => x"00", (0 + 1301) => x"00", (0 + 1302) => x"00", (0 + 1303) => x"00", (0 + 1304) => x"00", (0 + 1305) => x"00", (0 + 1306) => x"00", (0 + 1307) => x"00", (0 + 1308) => x"00", (0 + 1309) => x"00", (0 + 1310) => x"00", (0 + 1311) => x"00", (0 + 1312) => x"00", (0 + 1313) => x"00", (0 + 1314) => x"00", (0 + 1315) => x"00", (0 + 1316) => x"00", (0 + 1317) => x"00", (0 + 1318) => x"00", (0 + 1319) => x"00", (0 + 1320) => x"00", (0 + 1321) => x"00", (0 + 1322) => x"00", (0 + 1323) => x"00", (0 + 1324) => x"00", (0 + 1325) => x"00", (0 + 1326) => x"00", (0 + 1327) => x"00", (0 + 1328) => x"00", (0 + 1329) => x"00", (0 + 1330) => x"00", (0 + 1331) => x"00", (0 + 1332) => x"00", (0 + 1333) => x"00", (0 + 1334) => x"00", (0 + 1335) => x"00", (0 + 1336) => x"00", (0 + 1337) => x"00", (0 + 1338) => x"00", (0 + 1339) => x"00", (0 + 1340) => x"00", (0 + 1341) => x"00", (0 + 1342) => x"00", (0 + 1343) => x"00", (0 + 1344) => x"00", (0 + 1345) => x"00", (0 + 1346) => x"00", (0 + 1347) => x"00", (0 + 1348) => x"00", (0 + 1349) => x"00", (0 + 1350) => x"00", (0 + 1351) => x"00", (0 + 1352) => x"00", (0 + 1353) => x"00", (0 + 1354) => x"00", (0 + 1355) => x"00", (0 + 1356) => x"00", (0 + 1357) => x"00", (0 + 1358) => x"00", (0 + 1359) => x"00", (0 + 1360) => x"00", (0 + 1361) => x"00", (0 + 1362) => x"00", (0 + 1363) => x"00", (0 + 1364) => x"00", (0 + 1365) => x"00", (0 + 1366) => x"00", (0 + 1367) => x"00", (0 + 1368) => x"00", (0 + 1369) => x"00", (0 + 1370) => x"00", (0 + 1371) => x"00", (0 + 1372) => x"00", (0 + 1373) => x"00", (0 + 1374) => x"00", (0 + 1375) => x"00", (0 + 1376) => x"00", (0 + 1377) => x"00", (0 + 1378) => x"00", (0 + 1379) => x"00", (0 + 1380) => x"00", (0 + 1381) => x"00", (0 + 1382) => x"00", (0 + 1383) => x"00", (0 + 1384) => x"00", (0 + 1385) => x"00", (0 + 1386) => x"00", (0 + 1387) => x"00", (0 + 1388) => x"00", (0 + 1389) => x"00", (0 + 1390) => x"00", (0 + 1391) => x"00", (0 + 1392) => x"00", (0 + 1393) => x"00", (0 + 1394) => x"00", (0 + 1395) => x"00", (0 + 1396) => x"00", (0 + 1397) => x"00", (0 + 1398) => x"00", (0 + 1399) => x"00", (0 + 1400) => x"00", (0 + 1401) => x"00", (0 + 1402) => x"00", (0 + 1403) => x"00", (0 + 1404) => x"00", (0 + 1405) => x"00", (0 + 1406) => x"00", (0 + 1407) => x"00", (0 + 1408) => x"00", (0 + 1409) => x"00", (0 + 1410) => x"00", (0 + 1411) => x"00", (0 + 1412) => x"00", (0 + 1413) => x"00", (0 + 1414) => x"00", (0 + 1415) => x"00", (0 + 1416) => x"00", (0 + 1417) => x"00", (0 + 1418) => x"00", (0 + 1419) => x"00", (0 + 1420) => x"00", (0 + 1421) => x"00", (0 + 1422) => x"00", (0 + 1423) => x"00", (0 + 1424) => x"00", (0 + 1425) => x"00", (0 + 1426) => x"00", (0 + 1427) => x"00", (0 + 1428) => x"00", (0 + 1429) => x"00", (0 + 1430) => x"00", (0 + 1431) => x"00", (0 + 1432) => x"00", (0 + 1433) => x"00", (0 + 1434) => x"00", (0 + 1435) => x"00", (0 + 1436) => x"00", (0 + 1437) => x"00", (0 + 1438) => x"00", (0 + 1439) => x"00", (0 + 1440) => x"00", (0 + 1441) => x"00", (0 + 1442) => x"00", (0 + 1443) => x"00", (0 + 1444) => x"00", (0 + 1445) => x"00", (0 + 1446) => x"00", (0 + 1447) => x"00", (0 + 1448) => x"00", (0 + 1449) => x"00", (0 + 1450) => x"00", (0 + 1451) => x"00", (0 + 1452) => x"00", (0 + 1453) => x"00", (0 + 1454) => x"00", (0 + 1455) => x"00", (0 + 1456) => x"00", (0 + 1457) => x"00", (0 + 1458) => x"00", (0 + 1459) => x"00", (0 + 1460) => x"00", (0 + 1461) => x"00", (0 + 1462) => x"00", (0 + 1463) => x"00", (0 + 1464) => x"00", (0 + 1465) => x"00", (0 + 1466) => x"00", (0 + 1467) => x"00", (0 + 1468) => x"00", (0 + 1469) => x"00", (0 + 1470) => x"00", (0 + 1471) => x"00", (0 + 1472) => x"00", (0 + 1473) => x"00", (0 + 1474) => x"00", (0 + 1475) => x"00", (0 + 1476) => x"00", (0 + 1477) => x"00", (0 + 1478) => x"00", (0 + 1479) => x"00", (0 + 1480) => x"00", (0 + 1481) => x"00", (0 + 1482) => x"00", (0 + 1483) => x"00", (0 + 1484) => x"00", (0 + 1485) => x"00", (0 + 1486) => x"00", (0 + 1487) => x"00", (0 + 1488) => x"00", (0 + 1489) => x"00", (0 + 1490) => x"00", (0 + 1491) => x"00", (0 + 1492) => x"00", (0 + 1493) => x"00", (0 + 1494) => x"00", (0 + 1495) => x"00", (0 + 1496) => x"00", (0 + 1497) => x"00", (0 + 1498) => x"00", (0 + 1499) => x"00", (0 + 1500) => x"00", (0 + 1501) => x"00", (0 + 1502) => x"00", (0 + 1503) => x"00", (0 + 1504) => x"00", (0 + 1505) => x"00", (0 + 1506) => x"00", (0 + 1507) => x"00", (0 + 1508) => x"00", (0 + 1509) => x"00", (0 + 1510) => x"00", (0 + 1511) => x"00", (0 + 1512) => x"00", (0 + 1513) => x"00", (0 + 1514) => x"00", (0 + 1515) => x"00", (0 + 1516) => x"00", (0 + 1517) => x"00", (0 + 1518) => x"00", (0 + 1519) => x"00", (0 + 1520) => x"00", (0 + 1521) => x"00", (0 + 1522) => x"00", (0 + 1523) => x"00", (0 + 1524) => x"00", (0 + 1525) => x"00", (0 + 1526) => x"00", (0 + 1527) => x"00", (0 + 1528) => x"00", (0 + 1529) => x"00", (0 + 1530) => x"00", (0 + 1531) => x"00", (0 + 1532) => x"00", (0 + 1533) => x"00", (0 + 1534) => x"00", (0 + 1535) => x"00", (0 + 1536) => x"00", (0 + 1537) => x"00", (0 + 1538) => x"00", (0 + 1539) => x"00", (0 + 1540) => x"00", (0 + 1541) => x"00", (0 + 1542) => x"00", (0 + 1543) => x"00", (0 + 1544) => x"00", (0 + 1545) => x"00", (0 + 1546) => x"00", (0 + 1547) => x"00", (0 + 1548) => x"00", (0 + 1549) => x"00", (0 + 1550) => x"00", (0 + 1551) => x"00", (0 + 1552) => x"00", (0 + 1553) => x"00", (0 + 1554) => x"00", (0 + 1555) => x"00", (0 + 1556) => x"00", (0 + 1557) => x"00", (0 + 1558) => x"00", (0 + 1559) => x"00", (0 + 1560) => x"00", (0 + 1561) => x"00", (0 + 1562) => x"00", (0 + 1563) => x"00", (0 + 1564) => x"00", (0 + 1565) => x"00", (0 + 1566) => x"00", (0 + 1567) => x"00", (0 + 1568) => x"00", (0 + 1569) => x"00", (0 + 1570) => x"00", (0 + 1571) => x"00", (0 + 1572) => x"00", (0 + 1573) => x"00", (0 + 1574) => x"00", (0 + 1575) => x"00", (0 + 1576) => x"00", (0 + 1577) => x"00", (0 + 1578) => x"00", (0 + 1579) => x"00", (0 + 1580) => x"00", (0 + 1581) => x"00", (0 + 1582) => x"00", (0 + 1583) => x"00", (0 + 1584) => x"00", (0 + 1585) => x"00", (0 + 1586) => x"00", (0 + 1587) => x"00", (0 + 1588) => x"00", (0 + 1589) => x"00", (0 + 1590) => x"00", (0 + 1591) => x"00", (0 + 1592) => x"00", (0 + 1593) => x"00", (0 + 1594) => x"00", (0 + 1595) => x"00", (0 + 1596) => x"00", (0 + 1597) => x"00", (0 + 1598) => x"00", (0 + 1599) => x"00", (0 + 1600) => x"00", (0 + 1601) => x"00", (0 + 1602) => x"00", (0 + 1603) => x"00", (0 + 1604) => x"00", (0 + 1605) => x"00", (0 + 1606) => x"00", (0 + 1607) => x"00", (0 + 1608) => x"00", (0 + 1609) => x"00", (0 + 1610) => x"00", (0 + 1611) => x"00", (0 + 1612) => x"00", (0 + 1613) => x"00", (0 + 1614) => x"00", (0 + 1615) => x"00", (0 + 1616) => x"00", (0 + 1617) => x"00", (0 + 1618) => x"00", (0 + 1619) => x"00", (0 + 1620) => x"00", (0 + 1621) => x"00", (0 + 1622) => x"00", (0 + 1623) => x"00", (0 + 1624) => x"00", (0 + 1625) => x"00", (0 + 1626) => x"00", (0 + 1627) => x"00", (0 + 1628) => x"00", (0 + 1629) => x"00", (0 + 1630) => x"00", (0 + 1631) => x"00", (0 + 1632) => x"00", (0 + 1633) => x"00", (0 + 1634) => x"00", (0 + 1635) => x"00", (0 + 1636) => x"00", (0 + 1637) => x"00", (0 + 1638) => x"00", (0 + 1639) => x"00", (0 + 1640) => x"00", (0 + 1641) => x"00", (0 + 1642) => x"00", (0 + 1643) => x"00", (0 + 1644) => x"00", (0 + 1645) => x"00", (0 + 1646) => x"00", (0 + 1647) => x"00", (0 + 1648) => x"00", (0 + 1649) => x"00", (0 + 1650) => x"00", (0 + 1651) => x"00", (0 + 1652) => x"00", (0 + 1653) => x"00", (0 + 1654) => x"00", (0 + 1655) => x"00", (0 + 1656) => x"00", (0 + 1657) => x"00", (0 + 1658) => x"00", (0 + 1659) => x"00", (0 + 1660) => x"00", (0 + 1661) => x"00", (0 + 1662) => x"00", (0 + 1663) => x"00", (0 + 1664) => x"00", (0 + 1665) => x"00", (0 + 1666) => x"00", (0 + 1667) => x"00", (0 + 1668) => x"00", (0 + 1669) => x"00", (0 + 1670) => x"00", (0 + 1671) => x"00", (0 + 1672) => x"00", (0 + 1673) => x"00", (0 + 1674) => x"00", (0 + 1675) => x"00", (0 + 1676) => x"00", (0 + 1677) => x"00", (0 + 1678) => x"00", (0 + 1679) => x"00", (0 + 1680) => x"00", (0 + 1681) => x"00", (0 + 1682) => x"00", (0 + 1683) => x"00", (0 + 1684) => x"00", (0 + 1685) => x"00", (0 + 1686) => x"00", (0 + 1687) => x"00", (0 + 1688) => x"00", (0 + 1689) => x"00", (0 + 1690) => x"00", (0 + 1691) => x"00", (0 + 1692) => x"00", (0 + 1693) => x"00", (0 + 1694) => x"00", (0 + 1695) => x"00", (0 + 1696) => x"00", (0 + 1697) => x"00", (0 + 1698) => x"00", (0 + 1699) => x"00", (0 + 1700) => x"00", (0 + 1701) => x"00", (0 + 1702) => x"00", (0 + 1703) => x"00", (0 + 1704) => x"00", (0 + 1705) => x"00", (0 + 1706) => x"00", (0 + 1707) => x"00", (0 + 1708) => x"00", (0 + 1709) => x"00", (0 + 1710) => x"00", (0 + 1711) => x"00", (0 + 1712) => x"00", (0 + 1713) => x"00", (0 + 1714) => x"00", (0 + 1715) => x"00", (0 + 1716) => x"00", (0 + 1717) => x"00", (0 + 1718) => x"00", (0 + 1719) => x"00", (0 + 1720) => x"00", (0 + 1721) => x"00", (0 + 1722) => x"00", (0 + 1723) => x"00", (0 + 1724) => x"00", (0 + 1725) => x"00", (0 + 1726) => x"00", (0 + 1727) => x"00", (0 + 1728) => x"00", (0 + 1729) => x"00", (0 + 1730) => x"00", (0 + 1731) => x"00", (0 + 1732) => x"00", (0 + 1733) => x"00", (0 + 1734) => x"00", (0 + 1735) => x"00", (0 + 1736) => x"00", (0 + 1737) => x"00", (0 + 1738) => x"00", (0 + 1739) => x"00", (0 + 1740) => x"00", (0 + 1741) => x"00", (0 + 1742) => x"00", (0 + 1743) => x"00", (0 + 1744) => x"00", (0 + 1745) => x"00", (0 + 1746) => x"00", (0 + 1747) => x"00", (0 + 1748) => x"00", (0 + 1749) => x"00", (0 + 1750) => x"00", (0 + 1751) => x"00", (0 + 1752) => x"00", (0 + 1753) => x"00", (0 + 1754) => x"00", (0 + 1755) => x"00", (0 + 1756) => x"00", (0 + 1757) => x"00", (0 + 1758) => x"00", (0 + 1759) => x"00", (0 + 1760) => x"00", (0 + 1761) => x"00", (0 + 1762) => x"00", (0 + 1763) => x"00", (0 + 1764) => x"00", (0 + 1765) => x"00", (0 + 1766) => x"00", (0 + 1767) => x"00", (0 + 1768) => x"00", (0 + 1769) => x"00", (0 + 1770) => x"00", (0 + 1771) => x"00", (0 + 1772) => x"00", (0 + 1773) => x"00", (0 + 1774) => x"00", (0 + 1775) => x"00", (0 + 1776) => x"00", (0 + 1777) => x"00", (0 + 1778) => x"00", (0 + 1779) => x"00", (0 + 1780) => x"00", (0 + 1781) => x"00", (0 + 1782) => x"00", (0 + 1783) => x"00", (0 + 1784) => x"00", (0 + 1785) => x"00", (0 + 1786) => x"00", (0 + 1787) => x"00", (0 + 1788) => x"00", (0 + 1789) => x"00", (0 + 1790) => x"00", (0 + 1791) => x"00", (0 + 1792) => x"00", (0 + 1793) => x"00", (0 + 1794) => x"00", (0 + 1795) => x"00", (0 + 1796) => x"00", (0 + 1797) => x"00", (0 + 1798) => x"00", (0 + 1799) => x"00", (0 + 1800) => x"00", (0 + 1801) => x"00", (0 + 1802) => x"00", (0 + 1803) => x"00", (0 + 1804) => x"00", (0 + 1805) => x"00", (0 + 1806) => x"00", (0 + 1807) => x"00", (0 + 1808) => x"00", (0 + 1809) => x"00", (0 + 1810) => x"00", (0 + 1811) => x"00", (0 + 1812) => x"00", (0 + 1813) => x"00", (0 + 1814) => x"00", (0 + 1815) => x"00", (0 + 1816) => x"00", (0 + 1817) => x"00", (0 + 1818) => x"00", (0 + 1819) => x"00", (0 + 1820) => x"00", (0 + 1821) => x"00", (0 + 1822) => x"00", (0 + 1823) => x"00", (0 + 1824) => x"00", (0 + 1825) => x"00", (0 + 1826) => x"00", (0 + 1827) => x"00", (0 + 1828) => x"00", (0 + 1829) => x"00", (0 + 1830) => x"00", (0 + 1831) => x"00", (0 + 1832) => x"00", (0 + 1833) => x"00", (0 + 1834) => x"00", (0 + 1835) => x"00", (0 + 1836) => x"00", (0 + 1837) => x"00", (0 + 1838) => x"00", (0 + 1839) => x"00", (0 + 1840) => x"00", (0 + 1841) => x"00", (0 + 1842) => x"00", (0 + 1843) => x"00", (0 + 1844) => x"00", (0 + 1845) => x"00", (0 + 1846) => x"00", (0 + 1847) => x"00", (0 + 1848) => x"00", (0 + 1849) => x"00", (0 + 1850) => x"00", (0 + 1851) => x"00", (0 + 1852) => x"00", (0 + 1853) => x"00", (0 + 1854) => x"00", (0 + 1855) => x"00", (0 + 1856) => x"00", (0 + 1857) => x"00", (0 + 1858) => x"00", (0 + 1859) => x"00", (0 + 1860) => x"00", (0 + 1861) => x"00", (0 + 1862) => x"00", (0 + 1863) => x"00", (0 + 1864) => x"00", (0 + 1865) => x"00", (0 + 1866) => x"00", (0 + 1867) => x"00", (0 + 1868) => x"00", (0 + 1869) => x"00", (0 + 1870) => x"00", (0 + 1871) => x"00", (0 + 1872) => x"00", (0 + 1873) => x"00", (0 + 1874) => x"00", (0 + 1875) => x"00", (0 + 1876) => x"00", (0 + 1877) => x"00", (0 + 1878) => x"00", (0 + 1879) => x"00", (0 + 1880) => x"00", (0 + 1881) => x"00", (0 + 1882) => x"00", (0 + 1883) => x"00", (0 + 1884) => x"00", (0 + 1885) => x"00", (0 + 1886) => x"00", (0 + 1887) => x"00", (0 + 1888) => x"00", (0 + 1889) => x"00", (0 + 1890) => x"00", (0 + 1891) => x"00", (0 + 1892) => x"00", (0 + 1893) => x"00", (0 + 1894) => x"00", (0 + 1895) => x"00", (0 + 1896) => x"00", (0 + 1897) => x"00", (0 + 1898) => x"00", (0 + 1899) => x"00", (0 + 1900) => x"00", (0 + 1901) => x"00", (0 + 1902) => x"00", (0 + 1903) => x"00", (0 + 1904) => x"00", (0 + 1905) => x"00", (0 + 1906) => x"00", (0 + 1907) => x"00", (0 + 1908) => x"00", (0 + 1909) => x"00", (0 + 1910) => x"00", (0 + 1911) => x"00", (0 + 1912) => x"00", (0 + 1913) => x"00", (0 + 1914) => x"00", (0 + 1915) => x"00", (0 + 1916) => x"00", (0 + 1917) => x"00", (0 + 1918) => x"00", (0 + 1919) => x"00", (0 + 1920) => x"00", (0 + 1921) => x"00", (0 + 1922) => x"00", (0 + 1923) => x"00", (0 + 1924) => x"00", (0 + 1925) => x"00", (0 + 1926) => x"00", (0 + 1927) => x"00", (0 + 1928) => x"00", (0 + 1929) => x"00", (0 + 1930) => x"00", (0 + 1931) => x"00", (0 + 1932) => x"00", (0 + 1933) => x"00", (0 + 1934) => x"00", (0 + 1935) => x"00", (0 + 1936) => x"00", (0 + 1937) => x"00", (0 + 1938) => x"00", (0 + 1939) => x"00", (0 + 1940) => x"00", (0 + 1941) => x"00", (0 + 1942) => x"00", (0 + 1943) => x"00", (0 + 1944) => x"00", (0 + 1945) => x"00", (0 + 1946) => x"00", (0 + 1947) => x"00", (0 + 1948) => x"00", (0 + 1949) => x"00", (0 + 1950) => x"00", (0 + 1951) => x"00", (0 + 1952) => x"00", (0 + 1953) => x"00", (0 + 1954) => x"00", (0 + 1955) => x"00", (0 + 1956) => x"00", (0 + 1957) => x"00", (0 + 1958) => x"00", (0 + 1959) => x"00", (0 + 1960) => x"00", (0 + 1961) => x"00", (0 + 1962) => x"00", (0 + 1963) => x"00", (0 + 1964) => x"00", (0 + 1965) => x"00", (0 + 1966) => x"00", (0 + 1967) => x"00", (0 + 1968) => x"00", (0 + 1969) => x"00", (0 + 1970) => x"00", (0 + 1971) => x"00", (0 + 1972) => x"00", (0 + 1973) => x"00", (0 + 1974) => x"00", (0 + 1975) => x"00", (0 + 1976) => x"00", (0 + 1977) => x"00", (0 + 1978) => x"00", (0 + 1979) => x"00", (0 + 1980) => x"00", (0 + 1981) => x"00", (0 + 1982) => x"00", (0 + 1983) => x"00", (0 + 1984) => x"00", (0 + 1985) => x"00", (0 + 1986) => x"00", (0 + 1987) => x"00", (0 + 1988) => x"00", (0 + 1989) => x"00", (0 + 1990) => x"00", (0 + 1991) => x"00", (0 + 1992) => x"00", (0 + 1993) => x"00", (0 + 1994) => x"00", (0 + 1995) => x"00", (0 + 1996) => x"00", (0 + 1997) => x"00", (0 + 1998) => x"00", (0 + 1999) => x"00", (0 + 2000) => x"00", (0 + 2001) => x"00", (0 + 2002) => x"00", (0 + 2003) => x"00", (0 + 2004) => x"00", (0 + 2005) => x"00", (0 + 2006) => x"00", (0 + 2007) => x"00", (0 + 2008) => x"00", (0 + 2009) => x"00", (0 + 2010) => x"00", (0 + 2011) => x"00", (0 + 2012) => x"00", (0 + 2013) => x"00", (0 + 2014) => x"00", (0 + 2015) => x"00", (0 + 2016) => x"00", (0 + 2017) => x"00", (0 + 2018) => x"00", (0 + 2019) => x"00", (0 + 2020) => x"00", (0 + 2021) => x"00", (0 + 2022) => x"00", (0 + 2023) => x"00", (0 + 2024) => x"00", (0 + 2025) => x"00", (0 + 2026) => x"00", (0 + 2027) => x"00", (0 + 2028) => x"00", (0 + 2029) => x"00", (0 + 2030) => x"00", (0 + 2031) => x"00", (0 + 2032) => x"00", (0 + 2033) => x"00", (0 + 2034) => x"00", (0 + 2035) => x"00", (0 + 2036) => x"00", (0 + 2037) => x"00", (0 + 2038) => x"00", (0 + 2039) => x"00", (0 + 2040) => x"00", (0 + 2041) => x"00", (0 + 2042) => x"00", (0 + 2043) => x"00", (0 + 2044) => x"00", (0 + 2045) => x"00", (0 + 2046) => x"00", (0 + 2047) => x"00", (0 + 2048) => x"00", (0 + 2049) => x"00", (0 + 2050) => x"00", (0 + 2051) => x"00", (0 + 2052) => x"00", (0 + 2053) => x"00", (0 + 2054) => x"00", (0 + 2055) => x"00", (0 + 2056) => x"00", (0 + 2057) => x"00", (0 + 2058) => x"00", (0 + 2059) => x"00", (0 + 2060) => x"00", (0 + 2061) => x"00", (0 + 2062) => x"00", (0 + 2063) => x"00", (0 + 2064) => x"00", (0 + 2065) => x"00", (0 + 2066) => x"00", (0 + 2067) => x"00", (0 + 2068) => x"00", (0 + 2069) => x"00", (0 + 2070) => x"00", (0 + 2071) => x"00", (0 + 2072) => x"00", (0 + 2073) => x"00", (0 + 2074) => x"00", (0 + 2075) => x"00", (0 + 2076) => x"00", (0 + 2077) => x"00", (0 + 2078) => x"00", (0 + 2079) => x"00", (0 + 2080) => x"00", (0 + 2081) => x"00", (0 + 2082) => x"00", (0 + 2083) => x"00", (0 + 2084) => x"00", (0 + 2085) => x"00", (0 + 2086) => x"00", (0 + 2087) => x"00", (0 + 2088) => x"00", (0 + 2089) => x"00", (0 + 2090) => x"00", (0 + 2091) => x"00", (0 + 2092) => x"00", (0 + 2093) => x"00", (0 + 2094) => x"00", (0 + 2095) => x"00", (0 + 2096) => x"00", (0 + 2097) => x"00", (0 + 2098) => x"00", (0 + 2099) => x"00", (0 + 2100) => x"00", (0 + 2101) => x"00", (0 + 2102) => x"00", (0 + 2103) => x"00", (0 + 2104) => x"00", (0 + 2105) => x"00", (0 + 2106) => x"00", (0 + 2107) => x"00", (0 + 2108) => x"00", (0 + 2109) => x"00", (0 + 2110) => x"00", (0 + 2111) => x"00", (0 + 2112) => x"00", (0 + 2113) => x"00", (0 + 2114) => x"00", (0 + 2115) => x"00", (0 + 2116) => x"00", (0 + 2117) => x"00", (0 + 2118) => x"00", (0 + 2119) => x"00", (0 + 2120) => x"00", (0 + 2121) => x"00", (0 + 2122) => x"00", (0 + 2123) => x"00", (0 + 2124) => x"00", (0 + 2125) => x"00", (0 + 2126) => x"00", (0 + 2127) => x"00", (0 + 2128) => x"00", (0 + 2129) => x"00", (0 + 2130) => x"00", (0 + 2131) => x"00", (0 + 2132) => x"00", (0 + 2133) => x"00", (0 + 2134) => x"00", (0 + 2135) => x"00", (0 + 2136) => x"00", (0 + 2137) => x"00", (0 + 2138) => x"00", (0 + 2139) => x"00", (0 + 2140) => x"00", (0 + 2141) => x"00", (0 + 2142) => x"00", (0 + 2143) => x"00", (0 + 2144) => x"00", (0 + 2145) => x"00", (0 + 2146) => x"00", (0 + 2147) => x"00", (0 + 2148) => x"00", (0 + 2149) => x"00", (0 + 2150) => x"00", (0 + 2151) => x"00", (0 + 2152) => x"00", (0 + 2153) => x"00", (0 + 2154) => x"00", (0 + 2155) => x"00", (0 + 2156) => x"00", (0 + 2157) => x"00", (0 + 2158) => x"00", (0 + 2159) => x"00", (0 + 2160) => x"00", (0 + 2161) => x"00", (0 + 2162) => x"00", (0 + 2163) => x"00", (0 + 2164) => x"00", (0 + 2165) => x"00", (0 + 2166) => x"00", (0 + 2167) => x"00", (0 + 2168) => x"00", (0 + 2169) => x"00", (0 + 2170) => x"00", (0 + 2171) => x"00", (0 + 2172) => x"00", (0 + 2173) => x"00", (0 + 2174) => x"00", (0 + 2175) => x"00", (0 + 2176) => x"00", (0 + 2177) => x"00", (0 + 2178) => x"00", (0 + 2179) => x"00", (0 + 2180) => x"00", (0 + 2181) => x"00", (0 + 2182) => x"00", (0 + 2183) => x"00", (0 + 2184) => x"00", (0 + 2185) => x"00", (0 + 2186) => x"00", (0 + 2187) => x"00", (0 + 2188) => x"00", (0 + 2189) => x"00", (0 + 2190) => x"00", (0 + 2191) => x"00", (0 + 2192) => x"00", (0 + 2193) => x"00", (0 + 2194) => x"00", (0 + 2195) => x"00", (0 + 2196) => x"00", (0 + 2197) => x"00", (0 + 2198) => x"00", (0 + 2199) => x"00", (0 + 2200) => x"00", (0 + 2201) => x"00", (0 + 2202) => x"00", (0 + 2203) => x"00", (0 + 2204) => x"00", (0 + 2205) => x"00", (0 + 2206) => x"00", (0 + 2207) => x"00", (0 + 2208) => x"00", (0 + 2209) => x"00", (0 + 2210) => x"00", (0 + 2211) => x"00", (0 + 2212) => x"00", (0 + 2213) => x"00", (0 + 2214) => x"00", (0 + 2215) => x"00", (0 + 2216) => x"00", (0 + 2217) => x"00", (0 + 2218) => x"00", (0 + 2219) => x"00", (0 + 2220) => x"00", (0 + 2221) => x"00", (0 + 2222) => x"00", (0 + 2223) => x"00", (0 + 2224) => x"00", (0 + 2225) => x"00", (0 + 2226) => x"00", (0 + 2227) => x"00", (0 + 2228) => x"00", (0 + 2229) => x"00", (0 + 2230) => x"00", (0 + 2231) => x"00", (0 + 2232) => x"00", (0 + 2233) => x"00", (0 + 2234) => x"00", (0 + 2235) => x"00", (0 + 2236) => x"00", (0 + 2237) => x"00", (0 + 2238) => x"00", (0 + 2239) => x"00", (0 + 2240) => x"00", (0 + 2241) => x"00", (0 + 2242) => x"00", (0 + 2243) => x"00", (0 + 2244) => x"00", (0 + 2245) => x"00", (0 + 2246) => x"00", (0 + 2247) => x"00", (0 + 2248) => x"00", (0 + 2249) => x"00", (0 + 2250) => x"00", (0 + 2251) => x"00", (0 + 2252) => x"00", (0 + 2253) => x"00", (0 + 2254) => x"00", (0 + 2255) => x"00", (0 + 2256) => x"00", (0 + 2257) => x"00", (0 + 2258) => x"00", (0 + 2259) => x"00", (0 + 2260) => x"00", (0 + 2261) => x"00", (0 + 2262) => x"00", (0 + 2263) => x"00", (0 + 2264) => x"00", (0 + 2265) => x"00", (0 + 2266) => x"00", (0 + 2267) => x"00", (0 + 2268) => x"00", (0 + 2269) => x"00", (0 + 2270) => x"00", (0 + 2271) => x"00", (0 + 2272) => x"00", (0 + 2273) => x"00", (0 + 2274) => x"00", (0 + 2275) => x"00", (0 + 2276) => x"00", (0 + 2277) => x"00", (0 + 2278) => x"00", (0 + 2279) => x"00", (0 + 2280) => x"00", (0 + 2281) => x"00", (0 + 2282) => x"00", (0 + 2283) => x"00", (0 + 2284) => x"00", (0 + 2285) => x"00", (0 + 2286) => x"00", (0 + 2287) => x"00", (0 + 2288) => x"00", (0 + 2289) => x"00", (0 + 2290) => x"00", (0 + 2291) => x"00", (0 + 2292) => x"00", (0 + 2293) => x"00", (0 + 2294) => x"00", (0 + 2295) => x"00", (0 + 2296) => x"00", (0 + 2297) => x"00", (0 + 2298) => x"00", (0 + 2299) => x"00", (0 + 2300) => x"00", (0 + 2301) => x"00", (0 + 2302) => x"00", (0 + 2303) => x"00", (0 + 2304) => x"00", (0 + 2305) => x"00", (0 + 2306) => x"00", (0 + 2307) => x"00", (0 + 2308) => x"00", (0 + 2309) => x"00", (0 + 2310) => x"00", (0 + 2311) => x"00", (0 + 2312) => x"00", (0 + 2313) => x"00", (0 + 2314) => x"00", (0 + 2315) => x"00", (0 + 2316) => x"00", (0 + 2317) => x"00", (0 + 2318) => x"00", (0 + 2319) => x"00", (0 + 2320) => x"00", (0 + 2321) => x"00", (0 + 2322) => x"00", (0 + 2323) => x"00", (0 + 2324) => x"00", (0 + 2325) => x"00", (0 + 2326) => x"00", (0 + 2327) => x"00", (0 + 2328) => x"00", (0 + 2329) => x"00", (0 + 2330) => x"00", (0 + 2331) => x"00", (0 + 2332) => x"00", (0 + 2333) => x"00", (0 + 2334) => x"00", (0 + 2335) => x"00", (0 + 2336) => x"00", (0 + 2337) => x"00", (0 + 2338) => x"00", (0 + 2339) => x"00", (0 + 2340) => x"00", (0 + 2341) => x"00", (0 + 2342) => x"00", (0 + 2343) => x"00", (0 + 2344) => x"00", (0 + 2345) => x"00", (0 + 2346) => x"00", (0 + 2347) => x"00", (0 + 2348) => x"00", (0 + 2349) => x"00", (0 + 2350) => x"00", (0 + 2351) => x"00", (0 + 2352) => x"00", (0 + 2353) => x"00", (0 + 2354) => x"00", (0 + 2355) => x"00", (0 + 2356) => x"00", (0 + 2357) => x"00", (0 + 2358) => x"00", (0 + 2359) => x"00", (0 + 2360) => x"00", (0 + 2361) => x"00", (0 + 2362) => x"00", (0 + 2363) => x"00", (0 + 2364) => x"00", (0 + 2365) => x"00", (0 + 2366) => x"00", (0 + 2367) => x"00", (0 + 2368) => x"00", (0 + 2369) => x"00", (0 + 2370) => x"00", (0 + 2371) => x"00", (0 + 2372) => x"00", (0 + 2373) => x"00", (0 + 2374) => x"00", (0 + 2375) => x"00", (0 + 2376) => x"00", (0 + 2377) => x"00", (0 + 2378) => x"00", (0 + 2379) => x"00", (0 + 2380) => x"00", (0 + 2381) => x"00", (0 + 2382) => x"00", (0 + 2383) => x"00", (0 + 2384) => x"00", (0 + 2385) => x"00", (0 + 2386) => x"00", (0 + 2387) => x"00", (0 + 2388) => x"00", (0 + 2389) => x"00", (0 + 2390) => x"00", (0 + 2391) => x"00", (0 + 2392) => x"00", (0 + 2393) => x"00", (0 + 2394) => x"00", (0 + 2395) => x"00", (0 + 2396) => x"00", (0 + 2397) => x"00", (0 + 2398) => x"00", (0 + 2399) => x"00", (0 + 2400) => x"00", (0 + 2401) => x"00", (0 + 2402) => x"00", (0 + 2403) => x"00", (0 + 2404) => x"00", (0 + 2405) => x"00", (0 + 2406) => x"00", (0 + 2407) => x"00", (0 + 2408) => x"00", (0 + 2409) => x"00", (0 + 2410) => x"00", (0 + 2411) => x"00", (0 + 2412) => x"00", (0 + 2413) => x"00", (0 + 2414) => x"00", (0 + 2415) => x"00", (0 + 2416) => x"00", (0 + 2417) => x"00", (0 + 2418) => x"00", (0 + 2419) => x"00", (0 + 2420) => x"00", (0 + 2421) => x"00", (0 + 2422) => x"00", (0 + 2423) => x"00", (0 + 2424) => x"00", (0 + 2425) => x"00", (0 + 2426) => x"00", (0 + 2427) => x"00", (0 + 2428) => x"00", (0 + 2429) => x"00", (0 + 2430) => x"00", (0 + 2431) => x"00", (0 + 2432) => x"00", (0 + 2433) => x"00", (0 + 2434) => x"00", (0 + 2435) => x"00", (0 + 2436) => x"00", (0 + 2437) => x"00", (0 + 2438) => x"00", (0 + 2439) => x"00", (0 + 2440) => x"00", (0 + 2441) => x"00", (0 + 2442) => x"00", (0 + 2443) => x"00", (0 + 2444) => x"00", (0 + 2445) => x"00", (0 + 2446) => x"00", (0 + 2447) => x"00", (0 + 2448) => x"00", (0 + 2449) => x"00", (0 + 2450) => x"00", (0 + 2451) => x"00", (0 + 2452) => x"00", (0 + 2453) => x"00", (0 + 2454) => x"00", (0 + 2455) => x"00", (0 + 2456) => x"00", (0 + 2457) => x"00", (0 + 2458) => x"00", (0 + 2459) => x"00", (0 + 2460) => x"00", (0 + 2461) => x"00", (0 + 2462) => x"00", (0 + 2463) => x"00", (0 + 2464) => x"00", (0 + 2465) => x"00", (0 + 2466) => x"00", (0 + 2467) => x"00", (0 + 2468) => x"00", (0 + 2469) => x"00", (0 + 2470) => x"00", (0 + 2471) => x"00", (0 + 2472) => x"00", (0 + 2473) => x"00", (0 + 2474) => x"00", (0 + 2475) => x"00", (0 + 2476) => x"00", (0 + 2477) => x"00", (0 + 2478) => x"00", (0 + 2479) => x"00", (0 + 2480) => x"00", (0 + 2481) => x"00", (0 + 2482) => x"00", (0 + 2483) => x"00", (0 + 2484) => x"00", (0 + 2485) => x"00", (0 + 2486) => x"00", (0 + 2487) => x"00", (0 + 2488) => x"00", (0 + 2489) => x"00", (0 + 2490) => x"00", (0 + 2491) => x"00", (0 + 2492) => x"00", (0 + 2493) => x"00", (0 + 2494) => x"00", (0 + 2495) => x"00", (0 + 2496) => x"00", (0 + 2497) => x"00", (0 + 2498) => x"00", (0 + 2499) => x"00", (0 + 2500) => x"00", (0 + 2501) => x"00", (0 + 2502) => x"00", (0 + 2503) => x"00", (0 + 2504) => x"00", (0 + 2505) => x"00", (0 + 2506) => x"00", (0 + 2507) => x"00", (0 + 2508) => x"00", (0 + 2509) => x"00", (0 + 2510) => x"00", (0 + 2511) => x"00", (0 + 2512) => x"00", (0 + 2513) => x"00", (0 + 2514) => x"00", (0 + 2515) => x"00", (0 + 2516) => x"00", (0 + 2517) => x"00", (0 + 2518) => x"00", (0 + 2519) => x"00", (0 + 2520) => x"00", (0 + 2521) => x"00", (0 + 2522) => x"00", (0 + 2523) => x"00", (0 + 2524) => x"00", (0 + 2525) => x"00", (0 + 2526) => x"00", (0 + 2527) => x"00", (0 + 2528) => x"00", (0 + 2529) => x"00", (0 + 2530) => x"00", (0 + 2531) => x"00", (0 + 2532) => x"00", (0 + 2533) => x"00", (0 + 2534) => x"00", (0 + 2535) => x"00", (0 + 2536) => x"00", (0 + 2537) => x"00", (0 + 2538) => x"00", (0 + 2539) => x"00", (0 + 2540) => x"00", (0 + 2541) => x"00", (0 + 2542) => x"00", (0 + 2543) => x"00", (0 + 2544) => x"00", (0 + 2545) => x"00", (0 + 2546) => x"00", (0 + 2547) => x"00", (0 + 2548) => x"00", (0 + 2549) => x"00", (0 + 2550) => x"00", (0 + 2551) => x"00", (0 + 2552) => x"00", (0 + 2553) => x"00", (0 + 2554) => x"00", (0 + 2555) => x"00", (0 + 2556) => x"00", (0 + 2557) => x"00", (0 + 2558) => x"00", (0 + 2559) => x"00", (0 + 2560) => x"00", (0 + 2561) => x"00", (0 + 2562) => x"00", (0 + 2563) => x"00", (0 + 2564) => x"00", (0 + 2565) => x"00", (0 + 2566) => x"00", (0 + 2567) => x"00", (0 + 2568) => x"00", (0 + 2569) => x"00", (0 + 2570) => x"00", (0 + 2571) => x"00", (0 + 2572) => x"00", (0 + 2573) => x"00", (0 + 2574) => x"00", (0 + 2575) => x"00", (0 + 2576) => x"00", (0 + 2577) => x"00", (0 + 2578) => x"00", (0 + 2579) => x"00", (0 + 2580) => x"00", (0 + 2581) => x"00", (0 + 2582) => x"00", (0 + 2583) => x"00", (0 + 2584) => x"00", (0 + 2585) => x"00", (0 + 2586) => x"00", (0 + 2587) => x"00", (0 + 2588) => x"00", (0 + 2589) => x"00", (0 + 2590) => x"00", (0 + 2591) => x"00", (0 + 2592) => x"00", (0 + 2593) => x"00", (0 + 2594) => x"00", (0 + 2595) => x"00", (0 + 2596) => x"00", (0 + 2597) => x"00", (0 + 2598) => x"00", (0 + 2599) => x"00", (0 + 2600) => x"00", (0 + 2601) => x"00", (0 + 2602) => x"00", (0 + 2603) => x"00", (0 + 2604) => x"00", (0 + 2605) => x"00", (0 + 2606) => x"00", (0 + 2607) => x"00", (0 + 2608) => x"00", (0 + 2609) => x"00", (0 + 2610) => x"00", (0 + 2611) => x"00", (0 + 2612) => x"00", (0 + 2613) => x"00", (0 + 2614) => x"00", (0 + 2615) => x"00", (0 + 2616) => x"00", (0 + 2617) => x"00", (0 + 2618) => x"00", (0 + 2619) => x"00", (0 + 2620) => x"00", (0 + 2621) => x"00", (0 + 2622) => x"00", (0 + 2623) => x"00", (0 + 2624) => x"00", (0 + 2625) => x"00", (0 + 2626) => x"00", (0 + 2627) => x"00", (0 + 2628) => x"00", (0 + 2629) => x"00", (0 + 2630) => x"00", (0 + 2631) => x"00", (0 + 2632) => x"00", (0 + 2633) => x"00", (0 + 2634) => x"00", (0 + 2635) => x"00", (0 + 2636) => x"00", (0 + 2637) => x"00", (0 + 2638) => x"00", (0 + 2639) => x"00", (0 + 2640) => x"00", (0 + 2641) => x"00", (0 + 2642) => x"00", (0 + 2643) => x"00", (0 + 2644) => x"00", (0 + 2645) => x"00", (0 + 2646) => x"00", (0 + 2647) => x"00", (0 + 2648) => x"00", (0 + 2649) => x"00", (0 + 2650) => x"00", (0 + 2651) => x"00", (0 + 2652) => x"00", (0 + 2653) => x"00", (0 + 2654) => x"00", (0 + 2655) => x"00", (0 + 2656) => x"00", (0 + 2657) => x"00", (0 + 2658) => x"00", (0 + 2659) => x"00", (0 + 2660) => x"00", (0 + 2661) => x"00", (0 + 2662) => x"00", (0 + 2663) => x"00", (0 + 2664) => x"00", (0 + 2665) => x"00", (0 + 2666) => x"00", (0 + 2667) => x"00", (0 + 2668) => x"00", (0 + 2669) => x"00", (0 + 2670) => x"00", (0 + 2671) => x"00", (0 + 2672) => x"00", (0 + 2673) => x"00", (0 + 2674) => x"00", (0 + 2675) => x"00", (0 + 2676) => x"00", (0 + 2677) => x"00", (0 + 2678) => x"00", (0 + 2679) => x"00", (0 + 2680) => x"00", (0 + 2681) => x"00", (0 + 2682) => x"00", (0 + 2683) => x"00", (0 + 2684) => x"00", (0 + 2685) => x"00", (0 + 2686) => x"00", (0 + 2687) => x"00", (0 + 2688) => x"00", (0 + 2689) => x"00", (0 + 2690) => x"00", (0 + 2691) => x"00", (0 + 2692) => x"00", (0 + 2693) => x"00", (0 + 2694) => x"00", (0 + 2695) => x"00", (0 + 2696) => x"00", (0 + 2697) => x"00", (0 + 2698) => x"00", (0 + 2699) => x"00", (0 + 2700) => x"00", (0 + 2701) => x"00", (0 + 2702) => x"00", (0 + 2703) => x"00", (0 + 2704) => x"00", (0 + 2705) => x"00", (0 + 2706) => x"00", (0 + 2707) => x"00", (0 + 2708) => x"00", (0 + 2709) => x"00", (0 + 2710) => x"00", (0 + 2711) => x"00", (0 + 2712) => x"00", (0 + 2713) => x"00", (0 + 2714) => x"00", (0 + 2715) => x"00", (0 + 2716) => x"00", (0 + 2717) => x"00", (0 + 2718) => x"00", (0 + 2719) => x"00", (0 + 2720) => x"00", (0 + 2721) => x"00", (0 + 2722) => x"00", (0 + 2723) => x"00", (0 + 2724) => x"00", (0 + 2725) => x"00", (0 + 2726) => x"00", (0 + 2727) => x"00", (0 + 2728) => x"00", (0 + 2729) => x"00", (0 + 2730) => x"00", (0 + 2731) => x"00", (0 + 2732) => x"00", (0 + 2733) => x"00", (0 + 2734) => x"00", (0 + 2735) => x"00", (0 + 2736) => x"00", (0 + 2737) => x"00", (0 + 2738) => x"00", (0 + 2739) => x"00", (0 + 2740) => x"00", (0 + 2741) => x"00", (0 + 2742) => x"00", (0 + 2743) => x"00", (0 + 2744) => x"00", (0 + 2745) => x"00", (0 + 2746) => x"00", (0 + 2747) => x"00", (0 + 2748) => x"00", (0 + 2749) => x"00", (0 + 2750) => x"00", (0 + 2751) => x"00", (0 + 2752) => x"00", (0 + 2753) => x"00", (0 + 2754) => x"00", (0 + 2755) => x"00", (0 + 2756) => x"00", (0 + 2757) => x"00", (0 + 2758) => x"00", (0 + 2759) => x"00", (0 + 2760) => x"00", (0 + 2761) => x"00", (0 + 2762) => x"00", (0 + 2763) => x"00", (0 + 2764) => x"00", (0 + 2765) => x"00", (0 + 2766) => x"00", (0 + 2767) => x"00", (0 + 2768) => x"00", (0 + 2769) => x"00", (0 + 2770) => x"00", (0 + 2771) => x"00", (0 + 2772) => x"00", (0 + 2773) => x"00", (0 + 2774) => x"00", (0 + 2775) => x"00", (0 + 2776) => x"00", (0 + 2777) => x"00", (0 + 2778) => x"00", (0 + 2779) => x"00", (0 + 2780) => x"00", (0 + 2781) => x"00", (0 + 2782) => x"00", (0 + 2783) => x"00", (0 + 2784) => x"00", (0 + 2785) => x"00", (0 + 2786) => x"00", (0 + 2787) => x"00", (0 + 2788) => x"00", (0 + 2789) => x"00", (0 + 2790) => x"00", (0 + 2791) => x"00", (0 + 2792) => x"00", (0 + 2793) => x"00", (0 + 2794) => x"00", (0 + 2795) => x"00", (0 + 2796) => x"00", (0 + 2797) => x"00", (0 + 2798) => x"00", (0 + 2799) => x"00", (0 + 2800) => x"00", (0 + 2801) => x"00", (0 + 2802) => x"00", (0 + 2803) => x"00", (0 + 2804) => x"00", (0 + 2805) => x"00", (0 + 2806) => x"00", (0 + 2807) => x"00", (0 + 2808) => x"00", (0 + 2809) => x"00", (0 + 2810) => x"00", (0 + 2811) => x"00", (0 + 2812) => x"00", (0 + 2813) => x"00", (0 + 2814) => x"00", (0 + 2815) => x"00", (0 + 2816) => x"00", (0 + 2817) => x"00", (0 + 2818) => x"00", (0 + 2819) => x"00", (0 + 2820) => x"00", (0 + 2821) => x"00", (0 + 2822) => x"00", (0 + 2823) => x"00", (0 + 2824) => x"00", (0 + 2825) => x"00", (0 + 2826) => x"00", (0 + 2827) => x"00", (0 + 2828) => x"00", (0 + 2829) => x"00", (0 + 2830) => x"00", (0 + 2831) => x"00", (0 + 2832) => x"00", (0 + 2833) => x"00", (0 + 2834) => x"00", (0 + 2835) => x"00", (0 + 2836) => x"00", (0 + 2837) => x"00", (0 + 2838) => x"00", (0 + 2839) => x"00", (0 + 2840) => x"00", (0 + 2841) => x"00", (0 + 2842) => x"00", (0 + 2843) => x"00", (0 + 2844) => x"00", (0 + 2845) => x"00", (0 + 2846) => x"00", (0 + 2847) => x"00", (0 + 2848) => x"00", (0 + 2849) => x"00", (0 + 2850) => x"00", (0 + 2851) => x"00", (0 + 2852) => x"00", (0 + 2853) => x"00", (0 + 2854) => x"00", (0 + 2855) => x"00", (0 + 2856) => x"00", (0 + 2857) => x"00", (0 + 2858) => x"00", (0 + 2859) => x"00", (0 + 2860) => x"00", (0 + 2861) => x"00", (0 + 2862) => x"00", (0 + 2863) => x"00", (0 + 2864) => x"00", (0 + 2865) => x"00", (0 + 2866) => x"00", (0 + 2867) => x"00", (0 + 2868) => x"00", (0 + 2869) => x"00", (0 + 2870) => x"00", (0 + 2871) => x"00", (0 + 2872) => x"00", (0 + 2873) => x"00", (0 + 2874) => x"00", (0 + 2875) => x"00", (0 + 2876) => x"00", (0 + 2877) => x"00", (0 + 2878) => x"00", (0 + 2879) => x"00", (0 + 2880) => x"00", (0 + 2881) => x"00", (0 + 2882) => x"00", (0 + 2883) => x"00", (0 + 2884) => x"00", (0 + 2885) => x"00", (0 + 2886) => x"00", (0 + 2887) => x"00", (0 + 2888) => x"00", (0 + 2889) => x"00", (0 + 2890) => x"00", (0 + 2891) => x"00", (0 + 2892) => x"00", (0 + 2893) => x"00", (0 + 2894) => x"00", (0 + 2895) => x"00", (0 + 2896) => x"00", (0 + 2897) => x"00", (0 + 2898) => x"00", (0 + 2899) => x"00", (0 + 2900) => x"00", (0 + 2901) => x"00", (0 + 2902) => x"00", (0 + 2903) => x"00", (0 + 2904) => x"00", (0 + 2905) => x"00", (0 + 2906) => x"00", (0 + 2907) => x"00", (0 + 2908) => x"00", (0 + 2909) => x"00", (0 + 2910) => x"00", (0 + 2911) => x"00", (0 + 2912) => x"00", (0 + 2913) => x"00", (0 + 2914) => x"00", (0 + 2915) => x"00", (0 + 2916) => x"00", (0 + 2917) => x"00", (0 + 2918) => x"00", (0 + 2919) => x"00", (0 + 2920) => x"00", (0 + 2921) => x"00", (0 + 2922) => x"00", (0 + 2923) => x"00", (0 + 2924) => x"00", (0 + 2925) => x"00", (0 + 2926) => x"00", (0 + 2927) => x"00", (0 + 2928) => x"00", (0 + 2929) => x"00", (0 + 2930) => x"00", (0 + 2931) => x"00", (0 + 2932) => x"00", (0 + 2933) => x"00", (0 + 2934) => x"00", (0 + 2935) => x"00", (0 + 2936) => x"00", (0 + 2937) => x"00", (0 + 2938) => x"00", (0 + 2939) => x"00", (0 + 2940) => x"00", (0 + 2941) => x"00", (0 + 2942) => x"00", (0 + 2943) => x"00", (0 + 2944) => x"00", (0 + 2945) => x"00", (0 + 2946) => x"00", (0 + 2947) => x"00", (0 + 2948) => x"00", (0 + 2949) => x"00", (0 + 2950) => x"00", (0 + 2951) => x"00", (0 + 2952) => x"00", (0 + 2953) => x"00", (0 + 2954) => x"00", (0 + 2955) => x"00", (0 + 2956) => x"00", (0 + 2957) => x"00", (0 + 2958) => x"00", (0 + 2959) => x"00", (0 + 2960) => x"00", (0 + 2961) => x"00", (0 + 2962) => x"00", (0 + 2963) => x"00", (0 + 2964) => x"00", (0 + 2965) => x"00", (0 + 2966) => x"00", (0 + 2967) => x"00", (0 + 2968) => x"00", (0 + 2969) => x"00", (0 + 2970) => x"00", (0 + 2971) => x"00", (0 + 2972) => x"00", (0 + 2973) => x"00", (0 + 2974) => x"00", (0 + 2975) => x"00", (0 + 2976) => x"00", (0 + 2977) => x"00", (0 + 2978) => x"00", (0 + 2979) => x"00", (0 + 2980) => x"00", (0 + 2981) => x"00", (0 + 2982) => x"00", (0 + 2983) => x"00", (0 + 2984) => x"00", (0 + 2985) => x"00", (0 + 2986) => x"00", (0 + 2987) => x"00", (0 + 2988) => x"00", (0 + 2989) => x"00", (0 + 2990) => x"00", (0 + 2991) => x"00", (0 + 2992) => x"00", (0 + 2993) => x"00", (0 + 2994) => x"00", (0 + 2995) => x"00", (0 + 2996) => x"00", (0 + 2997) => x"00", (0 + 2998) => x"00", (0 + 2999) => x"00", (0 + 3000) => x"00", (0 + 3001) => x"00", (0 + 3002) => x"00", (0 + 3003) => x"00", (0 + 3004) => x"00", (0 + 3005) => x"00", (0 + 3006) => x"00", (0 + 3007) => x"00", (0 + 3008) => x"00", (0 + 3009) => x"00", (0 + 3010) => x"00", (0 + 3011) => x"00", (0 + 3012) => x"00", (0 + 3013) => x"00", (0 + 3014) => x"00", (0 + 3015) => x"00", (0 + 3016) => x"00", (0 + 3017) => x"00", (0 + 3018) => x"00", (0 + 3019) => x"00", (0 + 3020) => x"00", (0 + 3021) => x"00", (0 + 3022) => x"00", (0 + 3023) => x"00", (0 + 3024) => x"00", (0 + 3025) => x"00", (0 + 3026) => x"00", (0 + 3027) => x"00", (0 + 3028) => x"00", (0 + 3029) => x"00", (0 + 3030) => x"00", (0 + 3031) => x"00", (0 + 3032) => x"00", (0 + 3033) => x"00", (0 + 3034) => x"00", (0 + 3035) => x"00", (0 + 3036) => x"00", (0 + 3037) => x"00", (0 + 3038) => x"00", (0 + 3039) => x"00", (0 + 3040) => x"00", (0 + 3041) => x"00", (0 + 3042) => x"00", (0 + 3043) => x"00", (0 + 3044) => x"00", (0 + 3045) => x"00", (0 + 3046) => x"00", (0 + 3047) => x"00", (0 + 3048) => x"00", (0 + 3049) => x"00", (0 + 3050) => x"00", (0 + 3051) => x"00", (0 + 3052) => x"00", (0 + 3053) => x"00", (0 + 3054) => x"00", (0 + 3055) => x"00", (0 + 3056) => x"00", (0 + 3057) => x"00", (0 + 3058) => x"00", (0 + 3059) => x"00", (0 + 3060) => x"00", (0 + 3061) => x"00", (0 + 3062) => x"00", (0 + 3063) => x"00", (0 + 3064) => x"00", (0 + 3065) => x"00", (0 + 3066) => x"00", (0 + 3067) => x"00", (0 + 3068) => x"00", (0 + 3069) => x"00", (0 + 3070) => x"00", (0 + 3071) => x"00", (0 + 3072) => x"00", (0 + 3073) => x"00", (0 + 3074) => x"00", (0 + 3075) => x"00", (0 + 3076) => x"00", (0 + 3077) => x"00", (0 + 3078) => x"00", (0 + 3079) => x"00", (0 + 3080) => x"00", (0 + 3081) => x"00", (0 + 3082) => x"00", (0 + 3083) => x"00", (0 + 3084) => x"00", (0 + 3085) => x"00", (0 + 3086) => x"00", (0 + 3087) => x"00", (0 + 3088) => x"00", (0 + 3089) => x"00", (0 + 3090) => x"00", (0 + 3091) => x"00", (0 + 3092) => x"00", (0 + 3093) => x"00", (0 + 3094) => x"00", (0 + 3095) => x"00", (0 + 3096) => x"00", (0 + 3097) => x"00", (0 + 3098) => x"00", (0 + 3099) => x"00", (0 + 3100) => x"00", (0 + 3101) => x"00", (0 + 3102) => x"00", (0 + 3103) => x"00", (0 + 3104) => x"00", (0 + 3105) => x"00", (0 + 3106) => x"00", (0 + 3107) => x"00", (0 + 3108) => x"00", (0 + 3109) => x"00", (0 + 3110) => x"00", (0 + 3111) => x"00", (0 + 3112) => x"00", (0 + 3113) => x"00", (0 + 3114) => x"00", (0 + 3115) => x"00", (0 + 3116) => x"00", (0 + 3117) => x"00", (0 + 3118) => x"00", (0 + 3119) => x"00", (0 + 3120) => x"00", (0 + 3121) => x"00", (0 + 3122) => x"00", (0 + 3123) => x"00", (0 + 3124) => x"00", (0 + 3125) => x"00", (0 + 3126) => x"00", (0 + 3127) => x"00", (0 + 3128) => x"00", (0 + 3129) => x"00", (0 + 3130) => x"00", (0 + 3131) => x"00", (0 + 3132) => x"00", (0 + 3133) => x"00", (0 + 3134) => x"00", (0 + 3135) => x"00", (0 + 3136) => x"00", (0 + 3137) => x"00", (0 + 3138) => x"00", (0 + 3139) => x"00", (0 + 3140) => x"00", (0 + 3141) => x"00", (0 + 3142) => x"00", (0 + 3143) => x"00", (0 + 3144) => x"00", (0 + 3145) => x"00", (0 + 3146) => x"00", (0 + 3147) => x"00", (0 + 3148) => x"00", (0 + 3149) => x"00", (0 + 3150) => x"00", (0 + 3151) => x"00", (0 + 3152) => x"00", (0 + 3153) => x"00", (0 + 3154) => x"00", (0 + 3155) => x"00", (0 + 3156) => x"00", (0 + 3157) => x"00", (0 + 3158) => x"00", (0 + 3159) => x"00", (0 + 3160) => x"00", (0 + 3161) => x"00", (0 + 3162) => x"00", (0 + 3163) => x"00", (0 + 3164) => x"00", (0 + 3165) => x"00", (0 + 3166) => x"00", (0 + 3167) => x"00", (0 + 3168) => x"00", (0 + 3169) => x"00", (0 + 3170) => x"00", (0 + 3171) => x"00", (0 + 3172) => x"00", (0 + 3173) => x"00", (0 + 3174) => x"00", (0 + 3175) => x"00", (0 + 3176) => x"00", (0 + 3177) => x"00", (0 + 3178) => x"00", (0 + 3179) => x"00", (0 + 3180) => x"00", (0 + 3181) => x"00", (0 + 3182) => x"00", (0 + 3183) => x"00", (0 + 3184) => x"00", (0 + 3185) => x"00", (0 + 3186) => x"00", (0 + 3187) => x"00", (0 + 3188) => x"00", (0 + 3189) => x"00", (0 + 3190) => x"00", (0 + 3191) => x"00", (0 + 3192) => x"00", (0 + 3193) => x"00", (0 + 3194) => x"00", (0 + 3195) => x"00", (0 + 3196) => x"00", (0 + 3197) => x"00", (0 + 3198) => x"00", (0 + 3199) => x"00", (0 + 3200) => x"00", (0 + 3201) => x"00", (0 + 3202) => x"00", (0 + 3203) => x"00", (0 + 3204) => x"00", (0 + 3205) => x"00", (0 + 3206) => x"00", (0 + 3207) => x"00", (0 + 3208) => x"00", (0 + 3209) => x"00", (0 + 3210) => x"00", (0 + 3211) => x"00", (0 + 3212) => x"00", (0 + 3213) => x"00", (0 + 3214) => x"00", (0 + 3215) => x"00", (0 + 3216) => x"00", (0 + 3217) => x"00", (0 + 3218) => x"00", (0 + 3219) => x"00", (0 + 3220) => x"00", (0 + 3221) => x"00", (0 + 3222) => x"00", (0 + 3223) => x"00", (0 + 3224) => x"00", (0 + 3225) => x"00", (0 + 3226) => x"00", (0 + 3227) => x"00", (0 + 3228) => x"00", (0 + 3229) => x"00", (0 + 3230) => x"00", (0 + 3231) => x"00", (0 + 3232) => x"00", (0 + 3233) => x"00", (0 + 3234) => x"00", (0 + 3235) => x"00", (0 + 3236) => x"00", (0 + 3237) => x"00", (0 + 3238) => x"00", (0 + 3239) => x"00", (0 + 3240) => x"00", (0 + 3241) => x"00", (0 + 3242) => x"00", (0 + 3243) => x"00", (0 + 3244) => x"00", (0 + 3245) => x"00", (0 + 3246) => x"00", (0 + 3247) => x"00", (0 + 3248) => x"00", (0 + 3249) => x"00", (0 + 3250) => x"00", (0 + 3251) => x"00", (0 + 3252) => x"00", (0 + 3253) => x"00", (0 + 3254) => x"00", (0 + 3255) => x"00", (0 + 3256) => x"00", (0 + 3257) => x"00", (0 + 3258) => x"00", (0 + 3259) => x"00", (0 + 3260) => x"00", (0 + 3261) => x"00", (0 + 3262) => x"00", (0 + 3263) => x"00", (0 + 3264) => x"00", (0 + 3265) => x"00", (0 + 3266) => x"00", (0 + 3267) => x"00", (0 + 3268) => x"00", (0 + 3269) => x"00", (0 + 3270) => x"00", (0 + 3271) => x"00", (0 + 3272) => x"00", (0 + 3273) => x"00", (0 + 3274) => x"00", (0 + 3275) => x"00", (0 + 3276) => x"00", (0 + 3277) => x"00", (0 + 3278) => x"00", (0 + 3279) => x"00", (0 + 3280) => x"00", (0 + 3281) => x"00", (0 + 3282) => x"00", (0 + 3283) => x"00", (0 + 3284) => x"00", (0 + 3285) => x"00", (0 + 3286) => x"00", (0 + 3287) => x"00", (0 + 3288) => x"00", (0 + 3289) => x"00", (0 + 3290) => x"00", (0 + 3291) => x"00", (0 + 3292) => x"00", (0 + 3293) => x"00", (0 + 3294) => x"00", (0 + 3295) => x"00", (0 + 3296) => x"00", (0 + 3297) => x"00", (0 + 3298) => x"00", (0 + 3299) => x"00", (0 + 3300) => x"00", (0 + 3301) => x"00", (0 + 3302) => x"00", (0 + 3303) => x"00", (0 + 3304) => x"00", (0 + 3305) => x"00", (0 + 3306) => x"00", (0 + 3307) => x"00", (0 + 3308) => x"00", (0 + 3309) => x"00", (0 + 3310) => x"00", (0 + 3311) => x"00", (0 + 3312) => x"00", (0 + 3313) => x"00", (0 + 3314) => x"00", (0 + 3315) => x"00", (0 + 3316) => x"00", (0 + 3317) => x"00", (0 + 3318) => x"00", (0 + 3319) => x"00", (0 + 3320) => x"00", (0 + 3321) => x"00", (0 + 3322) => x"00", (0 + 3323) => x"00", (0 + 3324) => x"00", (0 + 3325) => x"00", (0 + 3326) => x"00", (0 + 3327) => x"00", (0 + 3328) => x"00", (0 + 3329) => x"00", (0 + 3330) => x"00", (0 + 3331) => x"00", (0 + 3332) => x"00", (0 + 3333) => x"00", (0 + 3334) => x"00", (0 + 3335) => x"00", (0 + 3336) => x"00", (0 + 3337) => x"00", (0 + 3338) => x"00", (0 + 3339) => x"00", (0 + 3340) => x"00", (0 + 3341) => x"00", (0 + 3342) => x"00", (0 + 3343) => x"00", (0 + 3344) => x"00", (0 + 3345) => x"00", (0 + 3346) => x"00", (0 + 3347) => x"00", (0 + 3348) => x"00", (0 + 3349) => x"00", (0 + 3350) => x"00", (0 + 3351) => x"00", (0 + 3352) => x"00", (0 + 3353) => x"00", (0 + 3354) => x"00", (0 + 3355) => x"00", (0 + 3356) => x"00", (0 + 3357) => x"00", (0 + 3358) => x"00", (0 + 3359) => x"00", (0 + 3360) => x"00", (0 + 3361) => x"00", (0 + 3362) => x"00", (0 + 3363) => x"00", (0 + 3364) => x"00", (0 + 3365) => x"00", (0 + 3366) => x"00", (0 + 3367) => x"00", (0 + 3368) => x"00", (0 + 3369) => x"00", (0 + 3370) => x"00", (0 + 3371) => x"00", (0 + 3372) => x"00", (0 + 3373) => x"00", (0 + 3374) => x"00", (0 + 3375) => x"00", (0 + 3376) => x"00", (0 + 3377) => x"00", (0 + 3378) => x"00", (0 + 3379) => x"00", (0 + 3380) => x"00", (0 + 3381) => x"00", (0 + 3382) => x"00", (0 + 3383) => x"00", (0 + 3384) => x"00", (0 + 3385) => x"00", (0 + 3386) => x"00", (0 + 3387) => x"00", (0 + 3388) => x"00", (0 + 3389) => x"00", (0 + 3390) => x"00", (0 + 3391) => x"00", (0 + 3392) => x"00", (0 + 3393) => x"00", (0 + 3394) => x"00", (0 + 3395) => x"00", (0 + 3396) => x"00", (0 + 3397) => x"00", (0 + 3398) => x"00", (0 + 3399) => x"00", (0 + 3400) => x"00", (0 + 3401) => x"00", (0 + 3402) => x"00", (0 + 3403) => x"00", (0 + 3404) => x"00", (0 + 3405) => x"00", (0 + 3406) => x"00", (0 + 3407) => x"00", (0 + 3408) => x"00", (0 + 3409) => x"00", (0 + 3410) => x"00", (0 + 3411) => x"00", (0 + 3412) => x"00", (0 + 3413) => x"00", (0 + 3414) => x"00", (0 + 3415) => x"00", (0 + 3416) => x"00", (0 + 3417) => x"00", (0 + 3418) => x"00", (0 + 3419) => x"00", (0 + 3420) => x"00", (0 + 3421) => x"00", (0 + 3422) => x"00", (0 + 3423) => x"00", (0 + 3424) => x"00", (0 + 3425) => x"00", (0 + 3426) => x"00", (0 + 3427) => x"00", (0 + 3428) => x"00", (0 + 3429) => x"00", (0 + 3430) => x"00", (0 + 3431) => x"00", (0 + 3432) => x"00", (0 + 3433) => x"00", (0 + 3434) => x"00", (0 + 3435) => x"00", (0 + 3436) => x"00", (0 + 3437) => x"00", (0 + 3438) => x"00", (0 + 3439) => x"00", (0 + 3440) => x"00", (0 + 3441) => x"00", (0 + 3442) => x"00", (0 + 3443) => x"00", (0 + 3444) => x"00", (0 + 3445) => x"00", (0 + 3446) => x"00", (0 + 3447) => x"00", (0 + 3448) => x"00", (0 + 3449) => x"00", (0 + 3450) => x"00", (0 + 3451) => x"00", (0 + 3452) => x"00", (0 + 3453) => x"00", (0 + 3454) => x"00", (0 + 3455) => x"00", (0 + 3456) => x"00", (0 + 3457) => x"00", (0 + 3458) => x"00", (0 + 3459) => x"00", (0 + 3460) => x"00", (0 + 3461) => x"00", (0 + 3462) => x"00", (0 + 3463) => x"00", (0 + 3464) => x"00", (0 + 3465) => x"00", (0 + 3466) => x"00", (0 + 3467) => x"00", (0 + 3468) => x"00", (0 + 3469) => x"00", (0 + 3470) => x"00", (0 + 3471) => x"00", (0 + 3472) => x"00", (0 + 3473) => x"00", (0 + 3474) => x"00", (0 + 3475) => x"00", (0 + 3476) => x"00", (0 + 3477) => x"00", (0 + 3478) => x"00", (0 + 3479) => x"00", (0 + 3480) => x"00", (0 + 3481) => x"00", (0 + 3482) => x"00", (0 + 3483) => x"00", (0 + 3484) => x"00", (0 + 3485) => x"00", (0 + 3486) => x"00", (0 + 3487) => x"00", (0 + 3488) => x"00", (0 + 3489) => x"00", (0 + 3490) => x"00", (0 + 3491) => x"00", (0 + 3492) => x"00", (0 + 3493) => x"00", (0 + 3494) => x"00", (0 + 3495) => x"00", (0 + 3496) => x"00", (0 + 3497) => x"00", (0 + 3498) => x"00", (0 + 3499) => x"00", (0 + 3500) => x"00", (0 + 3501) => x"00", (0 + 3502) => x"00", (0 + 3503) => x"00", (0 + 3504) => x"00", (0 + 3505) => x"00", (0 + 3506) => x"00", (0 + 3507) => x"00", (0 + 3508) => x"00", (0 + 3509) => x"00", (0 + 3510) => x"00", (0 + 3511) => x"00", (0 + 3512) => x"00", (0 + 3513) => x"00", (0 + 3514) => x"00", (0 + 3515) => x"00", (0 + 3516) => x"00", (0 + 3517) => x"00", (0 + 3518) => x"00", (0 + 3519) => x"00", (0 + 3520) => x"00", (0 + 3521) => x"00", (0 + 3522) => x"00", (0 + 3523) => x"00", (0 + 3524) => x"00", (0 + 3525) => x"00", (0 + 3526) => x"00", (0 + 3527) => x"00", (0 + 3528) => x"00", (0 + 3529) => x"00", (0 + 3530) => x"00", (0 + 3531) => x"00", (0 + 3532) => x"00", (0 + 3533) => x"00", (0 + 3534) => x"00", (0 + 3535) => x"00", (0 + 3536) => x"00", (0 + 3537) => x"00", (0 + 3538) => x"00", (0 + 3539) => x"00", (0 + 3540) => x"00", (0 + 3541) => x"00", (0 + 3542) => x"00", (0 + 3543) => x"00", (0 + 3544) => x"00", (0 + 3545) => x"00", (0 + 3546) => x"00", (0 + 3547) => x"00", (0 + 3548) => x"00", (0 + 3549) => x"00", (0 + 3550) => x"00", (0 + 3551) => x"00", (0 + 3552) => x"00", (0 + 3553) => x"00", (0 + 3554) => x"00", (0 + 3555) => x"00", (0 + 3556) => x"00", (0 + 3557) => x"00", (0 + 3558) => x"00", (0 + 3559) => x"00", (0 + 3560) => x"00", (0 + 3561) => x"00", (0 + 3562) => x"00", (0 + 3563) => x"00", (0 + 3564) => x"00", (0 + 3565) => x"00", (0 + 3566) => x"00", (0 + 3567) => x"00", (0 + 3568) => x"00", (0 + 3569) => x"00", (0 + 3570) => x"00", (0 + 3571) => x"00", (0 + 3572) => x"00", (0 + 3573) => x"00", (0 + 3574) => x"00", (0 + 3575) => x"00", (0 + 3576) => x"00", (0 + 3577) => x"00", (0 + 3578) => x"00", (0 + 3579) => x"00", (0 + 3580) => x"00", (0 + 3581) => x"00", (0 + 3582) => x"00", (0 + 3583) => x"00", (0 + 3584) => x"00", (0 + 3585) => x"00", (0 + 3586) => x"00", (0 + 3587) => x"00", (0 + 3588) => x"00", (0 + 3589) => x"00", (0 + 3590) => x"00", (0 + 3591) => x"00", (0 + 3592) => x"00", (0 + 3593) => x"00", (0 + 3594) => x"00", (0 + 3595) => x"00", (0 + 3596) => x"00", (0 + 3597) => x"00", (0 + 3598) => x"00", (0 + 3599) => x"00", (0 + 3600) => x"00", (0 + 3601) => x"00", (0 + 3602) => x"00", (0 + 3603) => x"00", (0 + 3604) => x"00", (0 + 3605) => x"00", (0 + 3606) => x"00", (0 + 3607) => x"00", (0 + 3608) => x"00", (0 + 3609) => x"00", (0 + 3610) => x"00", (0 + 3611) => x"00", (0 + 3612) => x"00", (0 + 3613) => x"00", (0 + 3614) => x"00", (0 + 3615) => x"00", (0 + 3616) => x"00", (0 + 3617) => x"00", (0 + 3618) => x"00", (0 + 3619) => x"00", (0 + 3620) => x"00", (0 + 3621) => x"00", (0 + 3622) => x"00", (0 + 3623) => x"00", (0 + 3624) => x"00", (0 + 3625) => x"00", (0 + 3626) => x"00", (0 + 3627) => x"00", (0 + 3628) => x"00", (0 + 3629) => x"00", (0 + 3630) => x"00", (0 + 3631) => x"00", (0 + 3632) => x"00", (0 + 3633) => x"00", (0 + 3634) => x"00", (0 + 3635) => x"00", (0 + 3636) => x"00", (0 + 3637) => x"00", (0 + 3638) => x"00", (0 + 3639) => x"00", (0 + 3640) => x"00", (0 + 3641) => x"00", (0 + 3642) => x"00", (0 + 3643) => x"00", (0 + 3644) => x"00", (0 + 3645) => x"00", (0 + 3646) => x"00", (0 + 3647) => x"00", (0 + 3648) => x"00", (0 + 3649) => x"00", (0 + 3650) => x"00", (0 + 3651) => x"00", (0 + 3652) => x"00", (0 + 3653) => x"00", (0 + 3654) => x"00", (0 + 3655) => x"00", (0 + 3656) => x"00", (0 + 3657) => x"00", (0 + 3658) => x"00", (0 + 3659) => x"00", (0 + 3660) => x"00", (0 + 3661) => x"00", (0 + 3662) => x"00", (0 + 3663) => x"00", (0 + 3664) => x"00", (0 + 3665) => x"00", (0 + 3666) => x"00", (0 + 3667) => x"00", (0 + 3668) => x"00", (0 + 3669) => x"00", (0 + 3670) => x"00", (0 + 3671) => x"00", (0 + 3672) => x"00", (0 + 3673) => x"00", (0 + 3674) => x"00", (0 + 3675) => x"00", (0 + 3676) => x"00", (0 + 3677) => x"00", (0 + 3678) => x"00", (0 + 3679) => x"00", (0 + 3680) => x"00", (0 + 3681) => x"00", (0 + 3682) => x"00", (0 + 3683) => x"00", (0 + 3684) => x"00", (0 + 3685) => x"00", (0 + 3686) => x"00", (0 + 3687) => x"00", (0 + 3688) => x"00", (0 + 3689) => x"00", (0 + 3690) => x"00", (0 + 3691) => x"00", (0 + 3692) => x"00", (0 + 3693) => x"00", (0 + 3694) => x"00", (0 + 3695) => x"00", (0 + 3696) => x"00", (0 + 3697) => x"00", (0 + 3698) => x"00", (0 + 3699) => x"00", (0 + 3700) => x"00", (0 + 3701) => x"00", (0 + 3702) => x"00", (0 + 3703) => x"00", (0 + 3704) => x"00", (0 + 3705) => x"00", (0 + 3706) => x"00", (0 + 3707) => x"00", (0 + 3708) => x"00", (0 + 3709) => x"00", (0 + 3710) => x"00", (0 + 3711) => x"00", (0 + 3712) => x"00", (0 + 3713) => x"00", (0 + 3714) => x"00", (0 + 3715) => x"00", (0 + 3716) => x"00", (0 + 3717) => x"00", (0 + 3718) => x"00", (0 + 3719) => x"00", (0 + 3720) => x"00", (0 + 3721) => x"00", (0 + 3722) => x"00", (0 + 3723) => x"00", (0 + 3724) => x"00", (0 + 3725) => x"00", (0 + 3726) => x"00", (0 + 3727) => x"00", (0 + 3728) => x"00", (0 + 3729) => x"00", (0 + 3730) => x"00", (0 + 3731) => x"00", (0 + 3732) => x"00", (0 + 3733) => x"00", (0 + 3734) => x"00", (0 + 3735) => x"00", (0 + 3736) => x"00", (0 + 3737) => x"00", (0 + 3738) => x"00", (0 + 3739) => x"00", (0 + 3740) => x"00", (0 + 3741) => x"00", (0 + 3742) => x"00", (0 + 3743) => x"00", (0 + 3744) => x"00", (0 + 3745) => x"00", (0 + 3746) => x"00", (0 + 3747) => x"00", (0 + 3748) => x"00", (0 + 3749) => x"00", (0 + 3750) => x"00", (0 + 3751) => x"00", (0 + 3752) => x"00", (0 + 3753) => x"00", (0 + 3754) => x"00", (0 + 3755) => x"00", (0 + 3756) => x"00", (0 + 3757) => x"00", (0 + 3758) => x"00", (0 + 3759) => x"00", (0 + 3760) => x"00", (0 + 3761) => x"00", (0 + 3762) => x"00", (0 + 3763) => x"00", (0 + 3764) => x"00", (0 + 3765) => x"00", (0 + 3766) => x"00", (0 + 3767) => x"00", (0 + 3768) => x"00", (0 + 3769) => x"00", (0 + 3770) => x"00", (0 + 3771) => x"00", (0 + 3772) => x"00", (0 + 3773) => x"00", (0 + 3774) => x"00", (0 + 3775) => x"00", (0 + 3776) => x"00", (0 + 3777) => x"00", (0 + 3778) => x"00", (0 + 3779) => x"00", (0 + 3780) => x"00", (0 + 3781) => x"00", (0 + 3782) => x"00", (0 + 3783) => x"00", (0 + 3784) => x"00", (0 + 3785) => x"00", (0 + 3786) => x"00", (0 + 3787) => x"00", (0 + 3788) => x"00", (0 + 3789) => x"00", (0 + 3790) => x"00", (0 + 3791) => x"00", (0 + 3792) => x"00", (0 + 3793) => x"00", (0 + 3794) => x"00", (0 + 3795) => x"00", (0 + 3796) => x"00", (0 + 3797) => x"00", (0 + 3798) => x"00", (0 + 3799) => x"00", (0 + 3800) => x"00", (0 + 3801) => x"00", (0 + 3802) => x"00", (0 + 3803) => x"00", (0 + 3804) => x"00", (0 + 3805) => x"00", (0 + 3806) => x"00", (0 + 3807) => x"00", (0 + 3808) => x"00", (0 + 3809) => x"00", (0 + 3810) => x"00", (0 + 3811) => x"00", (0 + 3812) => x"00", (0 + 3813) => x"00", (0 + 3814) => x"00", (0 + 3815) => x"00", (0 + 3816) => x"00", (0 + 3817) => x"00", (0 + 3818) => x"00", (0 + 3819) => x"00", (0 + 3820) => x"00", (0 + 3821) => x"00", (0 + 3822) => x"00", (0 + 3823) => x"00", (0 + 3824) => x"00", (0 + 3825) => x"00", (0 + 3826) => x"00", (0 + 3827) => x"00", (0 + 3828) => x"00", (0 + 3829) => x"00", (0 + 3830) => x"00", (0 + 3831) => x"00", (0 + 3832) => x"00", (0 + 3833) => x"00", (0 + 3834) => x"00", (0 + 3835) => x"00", (0 + 3836) => x"00", (0 + 3837) => x"00", (0 + 3838) => x"00", (0 + 3839) => x"00", (0 + 3840) => x"00", (0 + 3841) => x"00", (0 + 3842) => x"00", (0 + 3843) => x"00", (0 + 3844) => x"00", (0 + 3845) => x"00", (0 + 3846) => x"00", (0 + 3847) => x"00", (0 + 3848) => x"00", (0 + 3849) => x"00", (0 + 3850) => x"00", (0 + 3851) => x"00", (0 + 3852) => x"00", (0 + 3853) => x"00", (0 + 3854) => x"00", (0 + 3855) => x"00", (0 + 3856) => x"00", (0 + 3857) => x"00", (0 + 3858) => x"00", (0 + 3859) => x"00", (0 + 3860) => x"00", (0 + 3861) => x"00", (0 + 3862) => x"00", (0 + 3863) => x"00", (0 + 3864) => x"00", (0 + 3865) => x"00", (0 + 3866) => x"00", (0 + 3867) => x"00", (0 + 3868) => x"00", (0 + 3869) => x"00", (0 + 3870) => x"00", (0 + 3871) => x"00", (0 + 3872) => x"00", (0 + 3873) => x"00", (0 + 3874) => x"00", (0 + 3875) => x"00", (0 + 3876) => x"00", (0 + 3877) => x"00", (0 + 3878) => x"00", (0 + 3879) => x"00", (0 + 3880) => x"00", (0 + 3881) => x"00", (0 + 3882) => x"00", (0 + 3883) => x"00", (0 + 3884) => x"00", (0 + 3885) => x"00", (0 + 3886) => x"00", (0 + 3887) => x"00", (0 + 3888) => x"00", (0 + 3889) => x"00", (0 + 3890) => x"00", (0 + 3891) => x"00", (0 + 3892) => x"00", (0 + 3893) => x"00", (0 + 3894) => x"00", (0 + 3895) => x"00", (0 + 3896) => x"00", (0 + 3897) => x"00", (0 + 3898) => x"00", (0 + 3899) => x"00", (0 + 3900) => x"00", (0 + 3901) => x"00", (0 + 3902) => x"00", (0 + 3903) => x"00", (0 + 3904) => x"00", (0 + 3905) => x"00", (0 + 3906) => x"00", (0 + 3907) => x"00", (0 + 3908) => x"00", (0 + 3909) => x"00", (0 + 3910) => x"00", (0 + 3911) => x"00", (0 + 3912) => x"00", (0 + 3913) => x"00", (0 + 3914) => x"00", (0 + 3915) => x"00", (0 + 3916) => x"00", (0 + 3917) => x"00", (0 + 3918) => x"00", (0 + 3919) => x"00", (0 + 3920) => x"00", (0 + 3921) => x"00", (0 + 3922) => x"00", (0 + 3923) => x"00", (0 + 3924) => x"00", (0 + 3925) => x"00", (0 + 3926) => x"00", (0 + 3927) => x"00", (0 + 3928) => x"00", (0 + 3929) => x"00", (0 + 3930) => x"00", (0 + 3931) => x"00", (0 + 3932) => x"00", (0 + 3933) => x"00", (0 + 3934) => x"00", (0 + 3935) => x"00", (0 + 3936) => x"00", (0 + 3937) => x"00", (0 + 3938) => x"00", (0 + 3939) => x"00", (0 + 3940) => x"00", (0 + 3941) => x"00", (0 + 3942) => x"00", (0 + 3943) => x"00", (0 + 3944) => x"00", (0 + 3945) => x"00", (0 + 3946) => x"00", (0 + 3947) => x"00", (0 + 3948) => x"00", (0 + 3949) => x"00", (0 + 3950) => x"00", (0 + 3951) => x"00", (0 + 3952) => x"00", (0 + 3953) => x"00", (0 + 3954) => x"00", (0 + 3955) => x"00", (0 + 3956) => x"00", (0 + 3957) => x"00", (0 + 3958) => x"00", (0 + 3959) => x"00", (0 + 3960) => x"00", (0 + 3961) => x"00", (0 + 3962) => x"00", (0 + 3963) => x"00", (0 + 3964) => x"00", (0 + 3965) => x"00", (0 + 3966) => x"00", (0 + 3967) => x"00", (0 + 3968) => x"00", (0 + 3969) => x"00", (0 + 3970) => x"00", (0 + 3971) => x"00", (0 + 3972) => x"00", (0 + 3973) => x"00", (0 + 3974) => x"00", (0 + 3975) => x"00", (0 + 3976) => x"00", (0 + 3977) => x"00", (0 + 3978) => x"00", (0 + 3979) => x"00", (0 + 3980) => x"00", (0 + 3981) => x"00", (0 + 3982) => x"00", (0 + 3983) => x"00", (0 + 3984) => x"00", (0 + 3985) => x"00", (0 + 3986) => x"00", (0 + 3987) => x"00", (0 + 3988) => x"00", (0 + 3989) => x"00", (0 + 3990) => x"00", (0 + 3991) => x"00", (0 + 3992) => x"00", (0 + 3993) => x"00", (0 + 3994) => x"00", (0 + 3995) => x"00", (0 + 3996) => x"00", (0 + 3997) => x"00", (0 + 3998) => x"00", (0 + 3999) => x"00", (0 + 4000) => x"00", (0 + 4001) => x"00", (0 + 4002) => x"00", (0 + 4003) => x"00", (0 + 4004) => x"00", (0 + 4005) => x"00", (0 + 4006) => x"00", (0 + 4007) => x"00", (0 + 4008) => x"00", (0 + 4009) => x"00", (0 + 4010) => x"00", (0 + 4011) => x"00", (0 + 4012) => x"00", (0 + 4013) => x"00", (0 + 4014) => x"00", (0 + 4015) => x"00", (0 + 4016) => x"00", (0 + 4017) => x"00", (0 + 4018) => x"00", (0 + 4019) => x"00", (0 + 4020) => x"00", (0 + 4021) => x"00", (0 + 4022) => x"00", (0 + 4023) => x"00", (0 + 4024) => x"00", (0 + 4025) => x"00", (0 + 4026) => x"00", (0 + 4027) => x"00", (0 + 4028) => x"00", (0 + 4029) => x"00", (0 + 4030) => x"00", (0 + 4031) => x"00", (0 + 4032) => x"00", (0 + 4033) => x"00", (0 + 4034) => x"00", (0 + 4035) => x"00", (0 + 4036) => x"00", (0 + 4037) => x"00", (0 + 4038) => x"00", (0 + 4039) => x"00", (0 + 4040) => x"00", (0 + 4041) => x"00", (0 + 4042) => x"00", (0 + 4043) => x"00", (0 + 4044) => x"00", (0 + 4045) => x"00", (0 + 4046) => x"00", (0 + 4047) => x"00", (0 + 4048) => x"00", (0 + 4049) => x"00", (0 + 4050) => x"00", (0 + 4051) => x"00", (0 + 4052) => x"00", (0 + 4053) => x"00", (0 + 4054) => x"00", (0 + 4055) => x"00", (0 + 4056) => x"00", (0 + 4057) => x"00", (0 + 4058) => x"00", (0 + 4059) => x"00", (0 + 4060) => x"00", (0 + 4061) => x"00", (0 + 4062) => x"00", (0 + 4063) => x"00", (0 + 4064) => x"00", (0 + 4065) => x"00", (0 + 4066) => x"00", (0 + 4067) => x"00", (0 + 4068) => x"00", (0 + 4069) => x"00", (0 + 4070) => x"00", (0 + 4071) => x"00", (0 + 4072) => x"00", (0 + 4073) => x"00", (0 + 4074) => x"00", (0 + 4075) => x"00", (0 + 4076) => x"00", (0 + 4077) => x"00", (0 + 4078) => x"00", (0 + 4079) => x"00", (0 + 4080) => x"00", (0 + 4081) => x"00", (0 + 4082) => x"00", (0 + 4083) => x"00", (0 + 4084) => x"00", (0 + 4085) => x"00", (0 + 4086) => x"00", (0 + 4087) => x"00", (0 + 4088) => x"00", (0 + 4089) => x"00", (0 + 4090) => x"00", (0 + 4091) => x"00", (0 + 4092) => x"00", (0 + 4093) => x"00", (0 + 4094) => x"00", (0 + 4095) => x"00", 


