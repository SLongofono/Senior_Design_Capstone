(0 + 0) => x"00001137", (0 + 1) => x"8071011b", (0 + 2) => x"01411113", (0 + 3) => x"1400006f", (0 + 4) => x"06054663", (0 + 5) => x"09801637", (0 + 6) => x"00900593", (0 + 7) => x"00a00813", (0 + 8) => x"00461613", (0 + 9) => x"00100893", (0 + 10) => x"00050713", (0 + 11) => x"04a5d463", (0 + 12) => x"00100793", (0 + 13) => x"0307473b", (0 + 14) => x"0027969b", (0 + 15) => x"00f687bb", (0 + 16) => x"0017979b", (0 + 17) => x"fee5c8e3", (0 + 18) => x"02e787bb", (0 + 19) => x"40f5053b", (0 + 20) => x"0307071b", (0 + 21) => x"0ff77713", (0 + 22) => x"00464783", (0 + 23) => x"0ff7f793", (0 + 24) => x"fe078ce3", (0 + 25) => x"00e601a3", (0 + 26) => x"011602a3", (0 + 27) => x"fa051ee3", (0 + 28) => x"00008067", (0 + 29) => x"00000513", (0 + 30) => x"fd9ff06f", (0 + 31) => x"09801737", (0 + 32) => x"00471713", (0 + 33) => x"00474783", (0 + 34) => x"0ff7f793", (0 + 35) => x"fe078ce3", (0 + 36) => x"02d00793", (0 + 37) => x"00f701a3", (0 + 38) => x"00100793", (0 + 39) => x"40a0053b", (0 + 40) => x"00f702a3", (0 + 41) => x"f71ff06f", (0 + 42) => x"fe010113", (0 + 43) => x"00113c23", (0 + 44) => x"00813823", (0 + 45) => x"00913423", (0 + 46) => x"01213023", (0 + 47) => x"04050863", (0 + 48) => x"00100793", (0 + 49) => x"00050413", (0 + 50) => x"06f50263", (0 + 51) => x"00000493", (0 + 52) => x"00100913", (0 + 53) => x"fff4051b", (0 + 54) => x"fd1ff0ef", (0 + 55) => x"ffe4041b", (0 + 56) => x"009504bb", (0 + 57) => x"00040663", (0 + 58) => x"ff2416e3", (0 + 59) => x"0014849b", (0 + 60) => x"01813083", (0 + 61) => x"01013403", (0 + 62) => x"00048513", (0 + 63) => x"00013903", (0 + 64) => x"00813483", (0 + 65) => x"02010113", (0 + 66) => x"00008067", (0 + 67) => x"01813083", (0 + 68) => x"01013403", (0 + 69) => x"00000493", (0 + 70) => x"00048513", (0 + 71) => x"00013903", (0 + 72) => x"00813483", (0 + 73) => x"02010113", (0 + 74) => x"00008067", (0 + 75) => x"01813083", (0 + 76) => x"01013403", (0 + 77) => x"00100493", (0 + 78) => x"00048513", (0 + 79) => x"00013903", (0 + 80) => x"00813483", (0 + 81) => x"02010113", (0 + 82) => x"00008067", (0 + 83) => x"fe010113", (0 + 84) => x"01300793", (0 + 85) => x"00006737", (0 + 86) => x"01b79793", (0 + 87) => x"a5a7071b", (0 + 88) => x"00113c23", (0 + 89) => x"00813823", (0 + 90) => x"00913423", (0 + 91) => x"01213023", (0 + 92) => x"00e79023", (0 + 93) => x"098017b7", (0 + 94) => x"00000697", (0 + 95) => x"35068693", (0 + 96) => x"02100713", (0 + 97) => x"00479793", (0 + 98) => x"00100593", (0 + 99) => x"0047c603", (0 + 100) => x"0ff67613", (0 + 101) => x"fe060ce3", (0 + 102) => x"00e781a3", (0 + 103) => x"00b782a3", (0 + 104) => x"00168693", (0 + 105) => x"0006c703", (0 + 106) => x"fe0712e3", (0 + 107) => x"09801437", (0 + 108) => x"00441413", (0 + 109) => x"00100713", (0 + 110) => x"00100813", (0 + 111) => x"00200893", (0 + 112) => x"00a00313", (0 + 113) => x"00900513", (0 + 114) => x"00000617", (0 + 115) => x"32060613", (0 + 116) => x"04900693", (0 + 117) => x"00444783", (0 + 118) => x"0ff7f793", (0 + 119) => x"fe078ce3", (0 + 120) => x"00d401a3", (0 + 121) => x"00e402a3", (0 + 122) => x"00160613", (0 + 123) => x"00064683", (0 + 124) => x"fe0692e3", (0 + 125) => x"00000493", (0 + 126) => x"00000e13", (0 + 127) => x"00144783", (0 + 128) => x"0ff7f793", (0 + 129) => x"fe078ce3", (0 + 130) => x"00044683", (0 + 131) => x"00e40123", (0 + 132) => x"0ff6f693", (0 + 133) => x"fd06879b", (0 + 134) => x"0ff7f613", (0 + 135) => x"000e1a63", (0 + 136) => x"0ac56463", (0 + 137) => x"009784bb", (0 + 138) => x"00100e13", (0 + 139) => x"fd1ff06f", (0 + 140) => x"070e0e63", (0 + 141) => x"fd1e14e3", (0 + 142) => x"1a668463", (0 + 143) => x"00000597", (0 + 144) => x"2f458593", (0 + 145) => x"04900613", (0 + 146) => x"00444783", (0 + 147) => x"0ff7f793", (0 + 148) => x"fe078ce3", (0 + 149) => x"00c401a3", (0 + 150) => x"00e402a3", (0 + 151) => x"00158593", (0 + 152) => x"0005c603", (0 + 153) => x"fe0612e3", (0 + 154) => x"00444783", (0 + 155) => x"0ff7f793", (0 + 156) => x"fe078ce3", (0 + 157) => x"00d401a3", (0 + 158) => x"00e402a3", (0 + 159) => x"00000617", (0 + 160) => x"2dc60613", (0 + 161) => x"07c00693", (0 + 162) => x"00444783", (0 + 163) => x"0ff7f793", (0 + 164) => x"fe078ce3", (0 + 165) => x"00d401a3", (0 + 166) => x"00e402a3", (0 + 167) => x"00160613", (0 + 168) => x"00064683", (0 + 169) => x"fe0692e3", (0 + 170) => x"f4dff06f", (0 + 171) => x"08c56863", (0 + 172) => x"0024969b", (0 + 173) => x"009684bb", (0 + 174) => x"0014949b", (0 + 175) => x"009784bb", (0 + 176) => x"00200e13", (0 + 177) => x"f39ff06f", (0 + 178) => x"0e668463", (0 + 179) => x"00000597", (0 + 180) => x"26458593", (0 + 181) => x"04900613", (0 + 182) => x"00444783", (0 + 183) => x"0ff7f793", (0 + 184) => x"fe078ce3", (0 + 185) => x"00c401a3", (0 + 186) => x"00e402a3", (0 + 187) => x"00158593", (0 + 188) => x"0005c603", (0 + 189) => x"fe0612e3", (0 + 190) => x"00444783", (0 + 191) => x"0ff7f793", (0 + 192) => x"fe078ce3", (0 + 193) => x"00d401a3", (0 + 194) => x"00e402a3", (0 + 195) => x"00000617", (0 + 196) => x"23c60613", (0 + 197) => x"07c00693", (0 + 198) => x"00444783", (0 + 199) => x"0ff7f793", (0 + 200) => x"fe078ce3", (0 + 201) => x"00d401a3", (0 + 202) => x"00e402a3", (0 + 203) => x"00160613", (0 + 204) => x"00064683", (0 + 205) => x"fe0692e3", (0 + 206) => x"ec5ff06f", (0 + 207) => x"0a668263", (0 + 208) => x"00000597", (0 + 209) => x"1f058593", (0 + 210) => x"04900613", (0 + 211) => x"00444783", (0 + 212) => x"0ff7f793", (0 + 213) => x"fe078ce3", (0 + 214) => x"00c401a3", (0 + 215) => x"00e402a3", (0 + 216) => x"00158593", (0 + 217) => x"0005c603", (0 + 218) => x"fe0612e3", (0 + 219) => x"00444783", (0 + 220) => x"0ff7f793", (0 + 221) => x"fe078ce3", (0 + 222) => x"00d401a3", (0 + 223) => x"00e402a3", (0 + 224) => x"00000617", (0 + 225) => x"1d860613", (0 + 226) => x"07c00693", (0 + 227) => x"00444783", (0 + 228) => x"0ff7f793", (0 + 229) => x"fe078ce3", (0 + 230) => x"00d401a3", (0 + 231) => x"00e402a3", (0 + 232) => x"00160613", (0 + 233) => x"00064683", (0 + 234) => x"fe0692e3", (0 + 235) => x"e49ff06f", (0 + 236) => x"00000617", (0 + 237) => x"14860613", (0 + 238) => x"04e00693", (0 + 239) => x"00444783", (0 + 240) => x"0ff7f793", (0 + 241) => x"fe078ce3", (0 + 242) => x"00d401a3", (0 + 243) => x"00e402a3", (0 + 244) => x"00160613", (0 + 245) => x"00064683", (0 + 246) => x"fe0692e3", (0 + 247) => x"dedff06f", (0 + 248) => x"00048513", (0 + 249) => x"00000097", (0 + 250) => x"cc4080e7", (0 + 251) => x"00050913", (0 + 252) => x"00000697", (0 + 253) => x"18868693", (0 + 254) => x"00a00713", (0 + 255) => x"00100613", (0 + 256) => x"00444783", (0 + 257) => x"0ff7f793", (0 + 258) => x"fe078ce3", (0 + 259) => x"00e401a3", (0 + 260) => x"00c402a3", (0 + 261) => x"00168693", (0 + 262) => x"0006c703", (0 + 263) => x"fe0712e3", (0 + 264) => x"00048513", (0 + 265) => x"bedff0ef", (0 + 266) => x"00000697", (0 + 267) => x"17068693", (0 + 268) => x"07c00713", (0 + 269) => x"00100613", (0 + 270) => x"00444783", (0 + 271) => x"0ff7f793", (0 + 272) => x"fe078ce3", (0 + 273) => x"00e401a3", (0 + 274) => x"00c402a3", (0 + 275) => x"00168693", (0 + 276) => x"0006c703", (0 + 277) => x"fe0712e3", (0 + 278) => x"00090513", (0 + 279) => x"bb5ff0ef", (0 + 280) => x"00000697", (0 + 281) => x"14068693", (0 + 282) => x"07c00713", (0 + 283) => x"00100613", (0 + 284) => x"00444783", (0 + 285) => x"0ff7f793", (0 + 286) => x"fe078ce3", (0 + 287) => x"00e401a3", (0 + 288) => x"00c402a3", (0 + 289) => x"00168693", (0 + 290) => x"0006c703", (0 + 291) => x"fe0712e3", (0 + 292) => x"00000697", (0 + 293) => x"11868693", (0 + 294) => x"04900713", (0 + 295) => x"00100613", (0 + 296) => x"00444783", (0 + 297) => x"0ff7f793", (0 + 298) => x"fe078ce3", (0 + 299) => x"00e401a3", (0 + 300) => x"00c402a3", (0 + 301) => x"00168693", (0 + 302) => x"0006c703", (0 + 303) => x"fe0712e3", (0 + 304) => x"cf5ff06f", (0 + 305) => x"00000000", (0 + 306) => x"46212121", (0 + 307) => x"4e4f4249", (0 + 308) => x"49434341", (0 + 309) => x"52455320", (0 + 310) => x"21524556", (0 + 311) => x"0a0a2121", (0 + 312) => x"00000000", (0 + 313) => x"00000000", (0 + 314) => x"75706e49", (0 + 315) => x"61562074", (0 + 316) => x"3a65756c", (0 + 317) => x"00203e0a", (0 + 318) => x"6576654e", (0 + 319) => x"6f672072", (0 + 320) => x"20322074", (0 + 321) => x"69676964", (0 + 322) => x"66207374", (0 + 323) => x"6f6c6c6f", (0 + 324) => x"20646577", (0 + 325) => x"61207962", (0 + 326) => x"77656e20", (0 + 327) => x"656e696c", (0 + 328) => x"7274202c", (0 + 329) => x"67612079", (0 + 330) => x"216e6961", (0 + 331) => x"000a0a21", (0 + 332) => x"61766e49", (0 + 333) => x"2064696c", (0 + 334) => x"72616843", (0 + 335) => x"65746361", (0 + 336) => x"007c2072", (0 + 337) => x"00000000", (0 + 338) => x"6b73207c", (0 + 339) => x"69707069", (0 + 340) => x"2121676e", (0 + 341) => x"00000a21", (0 + 342) => x"6769207c", (0 + 343) => x"69726f6e", (0 + 344) => x"7020676e", (0 + 345) => x"69766572", (0 + 346) => x"2073756f", (0 + 347) => x"756c6176", (0 + 348) => x"21217365", (0 + 349) => x"00000a21", (0 + 350) => x"6269660a", (0 + 351) => x"63616e6f", (0 + 352) => x"73206963", (0 + 353) => x"65757165", (0 + 354) => x"2065636e", (0 + 355) => x"7c207461", (0 + 356) => x"00000000", (0 + 357) => x"00000000", (0 + 358) => x"7369207c", (0 + 359) => x"00007c20", (0 + 360) => x"000a0a7c", (0 + 361) => x"00000000", (0 + 362) => x"75706e49", (0 + 363) => x"6e412074", (0 + 364) => x"6568746f", (0 + 365) => x"3f3f3f72", (0 + 366) => x"00000a3f", (0 + 367) => x"00000000", (0 + 368) => x"00000000", (0 + 369) => x"00000000", (0 + 370) => x"00000000", (0 + 371) => x"00000000", (0 + 372) => x"00000000", (0 + 373) => x"00000000", (0 + 374) => x"00000000", (0 + 375) => x"00000000", (0 + 376) => x"00000000", (0 + 377) => x"00000000", (0 + 378) => x"00000000", (0 + 379) => x"00000000", (0 + 380) => x"00000000", (0 + 381) => x"00000000", (0 + 382) => x"00000000", (0 + 383) => x"00000000", (0 + 384) => x"00000000", (0 + 385) => x"00000000", (0 + 386) => x"00000000", (0 + 387) => x"00000000", (0 + 388) => x"00000000", (0 + 389) => x"00000000", (0 + 390) => x"00000000", (0 + 391) => x"00000000", (0 + 392) => x"00000000", (0 + 393) => x"00000000", (0 + 394) => x"00000000", (0 + 395) => x"00000000", (0 + 396) => x"00000000", (0 + 397) => x"00000000", (0 + 398) => x"00000000", (0 + 399) => x"00000000", (0 + 400) => x"00000000", (0 + 401) => x"00000000", (0 + 402) => x"00000000", (0 + 403) => x"00000000", (0 + 404) => x"00000000", (0 + 405) => x"00000000", (0 + 406) => x"00000000", (0 + 407) => x"00000000", (0 + 408) => x"00000000", (0 + 409) => x"00000000", (0 + 410) => x"00000000", (0 + 411) => x"00000000", (0 + 412) => x"00000000", (0 + 413) => x"00000000", (0 + 414) => x"00000000", (0 + 415) => x"00000000", (0 + 416) => x"00000000", (0 + 417) => x"00000000", (0 + 418) => x"00000000", (0 + 419) => x"00000000", (0 + 420) => x"00000000", (0 + 421) => x"00000000", (0 + 422) => x"00000000", (0 + 423) => x"00000000", (0 + 424) => x"00000000", (0 + 425) => x"00000000", (0 + 426) => x"00000000", (0 + 427) => x"00000000", (0 + 428) => x"00000000", (0 + 429) => x"00000000", (0 + 430) => x"00000000", (0 + 431) => x"00000000", (0 + 432) => x"00000000", (0 + 433) => x"00000000", (0 + 434) => x"00000000", (0 + 435) => x"00000000", (0 + 436) => x"00000000", (0 + 437) => x"00000000", (0 + 438) => x"00000000", (0 + 439) => x"00000000", (0 + 440) => x"00000000", (0 + 441) => x"00000000", (0 + 442) => x"00000000", (0 + 443) => x"00000000", (0 + 444) => x"00000000", (0 + 445) => x"00000000", (0 + 446) => x"00000000", (0 + 447) => x"00000000", (0 + 448) => x"00000000", (0 + 449) => x"00000000", (0 + 450) => x"00000000", (0 + 451) => x"00000000", (0 + 452) => x"00000000", (0 + 453) => x"00000000", (0 + 454) => x"00000000", (0 + 455) => x"00000000", (0 + 456) => x"00000000", (0 + 457) => x"00000000", (0 + 458) => x"00000000", (0 + 459) => x"00000000", (0 + 460) => x"00000000", (0 + 461) => x"00000000", (0 + 462) => x"00000000", (0 + 463) => x"00000000", (0 + 464) => x"00000000", (0 + 465) => x"00000000", (0 + 466) => x"00000000", (0 + 467) => x"00000000", (0 + 468) => x"00000000", (0 + 469) => x"00000000", (0 + 470) => x"00000000", (0 + 471) => x"00000000", (0 + 472) => x"00000000", (0 + 473) => x"00000000", (0 + 474) => x"00000000", (0 + 475) => x"00000000", (0 + 476) => x"00000000", (0 + 477) => x"00000000", (0 + 478) => x"00000000", (0 + 479) => x"00000000", (0 + 480) => x"00000000", (0 + 481) => x"00000000", (0 + 482) => x"00000000", (0 + 483) => x"00000000", (0 + 484) => x"00000000", (0 + 485) => x"00000000", (0 + 486) => x"00000000", (0 + 487) => x"00000000", (0 + 488) => x"00000000", (0 + 489) => x"00000000", (0 + 490) => x"00000000", (0 + 491) => x"00000000", (0 + 492) => x"00000000", (0 + 493) => x"00000000", (0 + 494) => x"00000000", (0 + 495) => x"00000000", (0 + 496) => x"00000000", (0 + 497) => x"00000000", (0 + 498) => x"00000000", (0 + 499) => x"00000000", (0 + 500) => x"00000000", (0 + 501) => x"00000000", (0 + 502) => x"00000000", (0 + 503) => x"00000000", (0 + 504) => x"00000000", (0 + 505) => x"00000000", (0 + 506) => x"00000000", (0 + 507) => x"00000000", (0 + 508) => x"00000000", (0 + 509) => x"00000000", (0 + 510) => x"00000000", (0 + 511) => x"00000000", (0 + 512) => x"00000000", (0 + 513) => x"00000000", (0 + 514) => x"00000000", (0 + 515) => x"00000000", (0 + 516) => x"00000000", (0 + 517) => x"00000000", (0 + 518) => x"00000000", (0 + 519) => x"00000000", (0 + 520) => x"00000000", (0 + 521) => x"00000000", (0 + 522) => x"00000000", (0 + 523) => x"00000000", (0 + 524) => x"00000000", (0 + 525) => x"00000000", (0 + 526) => x"00000000", (0 + 527) => x"00000000", (0 + 528) => x"00000000", (0 + 529) => x"00000000", (0 + 530) => x"00000000", (0 + 531) => x"00000000", (0 + 532) => x"00000000", (0 + 533) => x"00000000", (0 + 534) => x"00000000", (0 + 535) => x"00000000", (0 + 536) => x"00000000", (0 + 537) => x"00000000", (0 + 538) => x"00000000", (0 + 539) => x"00000000", (0 + 540) => x"00000000", (0 + 541) => x"00000000", (0 + 542) => x"00000000", (0 + 543) => x"00000000", (0 + 544) => x"00000000", (0 + 545) => x"00000000", (0 + 546) => x"00000000", (0 + 547) => x"00000000", (0 + 548) => x"00000000", (0 + 549) => x"00000000", (0 + 550) => x"00000000", (0 + 551) => x"00000000", (0 + 552) => x"00000000", (0 + 553) => x"00000000", (0 + 554) => x"00000000", (0 + 555) => x"00000000", (0 + 556) => x"00000000", (0 + 557) => x"00000000", (0 + 558) => x"00000000", (0 + 559) => x"00000000", (0 + 560) => x"00000000", (0 + 561) => x"00000000", (0 + 562) => x"00000000", (0 + 563) => x"00000000", (0 + 564) => x"00000000", (0 + 565) => x"00000000", (0 + 566) => x"00000000", (0 + 567) => x"00000000", (0 + 568) => x"00000000", (0 + 569) => x"00000000", (0 + 570) => x"00000000", (0 + 571) => x"00000000", (0 + 572) => x"00000000", (0 + 573) => x"00000000", (0 + 574) => x"00000000", (0 + 575) => x"00000000", (0 + 576) => x"00000000", (0 + 577) => x"00000000", (0 + 578) => x"00000000", (0 + 579) => x"00000000", (0 + 580) => x"00000000", (0 + 581) => x"00000000", (0 + 582) => x"00000000", (0 + 583) => x"00000000", (0 + 584) => x"00000000", (0 + 585) => x"00000000", (0 + 586) => x"00000000", (0 + 587) => x"00000000", (0 + 588) => x"00000000", (0 + 589) => x"00000000", (0 + 590) => x"00000000", (0 + 591) => x"00000000", (0 + 592) => x"00000000", (0 + 593) => x"00000000", (0 + 594) => x"00000000", (0 + 595) => x"00000000", (0 + 596) => x"00000000", (0 + 597) => x"00000000", (0 + 598) => x"00000000", (0 + 599) => x"00000000", (0 + 600) => x"00000000", (0 + 601) => x"00000000", (0 + 602) => x"00000000", (0 + 603) => x"00000000", (0 + 604) => x"00000000", (0 + 605) => x"00000000", (0 + 606) => x"00000000", (0 + 607) => x"00000000", (0 + 608) => x"00000000", (0 + 609) => x"00000000", (0 + 610) => x"00000000", (0 + 611) => x"00000000", (0 + 612) => x"00000000", (0 + 613) => x"00000000", (0 + 614) => x"00000000", (0 + 615) => x"00000000", (0 + 616) => x"00000000", (0 + 617) => x"00000000", (0 + 618) => x"00000000", (0 + 619) => x"00000000", (0 + 620) => x"00000000", (0 + 621) => x"00000000", (0 + 622) => x"00000000", (0 + 623) => x"00000000", (0 + 624) => x"00000000", (0 + 625) => x"00000000", (0 + 626) => x"00000000", (0 + 627) => x"00000000", (0 + 628) => x"00000000", (0 + 629) => x"00000000", (0 + 630) => x"00000000", (0 + 631) => x"00000000", (0 + 632) => x"00000000", (0 + 633) => x"00000000", (0 + 634) => x"00000000", (0 + 635) => x"00000000", (0 + 636) => x"00000000", (0 + 637) => x"00000000", (0 + 638) => x"00000000", (0 + 639) => x"00000000", (0 + 640) => x"00000000", (0 + 641) => x"00000000", (0 + 642) => x"00000000", (0 + 643) => x"00000000", (0 + 644) => x"00000000", (0 + 645) => x"00000000", (0 + 646) => x"00000000", (0 + 647) => x"00000000", (0 + 648) => x"00000000", (0 + 649) => x"00000000", (0 + 650) => x"00000000", (0 + 651) => x"00000000", (0 + 652) => x"00000000", (0 + 653) => x"00000000", (0 + 654) => x"00000000", (0 + 655) => x"00000000", (0 + 656) => x"00000000", (0 + 657) => x"00000000", (0 + 658) => x"00000000", (0 + 659) => x"00000000", (0 + 660) => x"00000000", (0 + 661) => x"00000000", (0 + 662) => x"00000000", (0 + 663) => x"00000000", (0 + 664) => x"00000000", (0 + 665) => x"00000000", (0 + 666) => x"00000000", (0 + 667) => x"00000000", (0 + 668) => x"00000000", (0 + 669) => x"00000000", (0 + 670) => x"00000000", (0 + 671) => x"00000000", (0 + 672) => x"00000000", (0 + 673) => x"00000000", (0 + 674) => x"00000000", (0 + 675) => x"00000000", (0 + 676) => x"00000000", (0 + 677) => x"00000000", (0 + 678) => x"00000000", (0 + 679) => x"00000000", (0 + 680) => x"00000000", (0 + 681) => x"00000000", (0 + 682) => x"00000000", (0 + 683) => x"00000000", (0 + 684) => x"00000000", (0 + 685) => x"00000000", (0 + 686) => x"00000000", (0 + 687) => x"00000000", (0 + 688) => x"00000000", (0 + 689) => x"00000000", (0 + 690) => x"00000000", (0 + 691) => x"00000000", (0 + 692) => x"00000000", (0 + 693) => x"00000000", (0 + 694) => x"00000000", (0 + 695) => x"00000000", (0 + 696) => x"00000000", (0 + 697) => x"00000000", (0 + 698) => x"00000000", (0 + 699) => x"00000000", (0 + 700) => x"00000000", (0 + 701) => x"00000000", (0 + 702) => x"00000000", (0 + 703) => x"00000000", (0 + 704) => x"00000000", (0 + 705) => x"00000000", (0 + 706) => x"00000000", (0 + 707) => x"00000000", (0 + 708) => x"00000000", (0 + 709) => x"00000000", (0 + 710) => x"00000000", (0 + 711) => x"00000000", (0 + 712) => x"00000000", (0 + 713) => x"00000000", (0 + 714) => x"00000000", (0 + 715) => x"00000000", (0 + 716) => x"00000000", (0 + 717) => x"00000000", (0 + 718) => x"00000000", (0 + 719) => x"00000000", (0 + 720) => x"00000000", (0 + 721) => x"00000000", (0 + 722) => x"00000000", (0 + 723) => x"00000000", (0 + 724) => x"00000000", (0 + 725) => x"00000000", (0 + 726) => x"00000000", (0 + 727) => x"00000000", (0 + 728) => x"00000000", (0 + 729) => x"00000000", (0 + 730) => x"00000000", (0 + 731) => x"00000000", (0 + 732) => x"00000000", (0 + 733) => x"00000000", (0 + 734) => x"00000000", (0 + 735) => x"00000000", (0 + 736) => x"00000000", (0 + 737) => x"00000000", (0 + 738) => x"00000000", (0 + 739) => x"00000000", (0 + 740) => x"00000000", (0 + 741) => x"00000000", (0 + 742) => x"00000000", (0 + 743) => x"00000000", (0 + 744) => x"00000000", (0 + 745) => x"00000000", (0 + 746) => x"00000000", (0 + 747) => x"00000000", (0 + 748) => x"00000000", (0 + 749) => x"00000000", (0 + 750) => x"00000000", (0 + 751) => x"00000000", (0 + 752) => x"00000000", (0 + 753) => x"00000000", (0 + 754) => x"00000000", (0 + 755) => x"00000000", (0 + 756) => x"00000000", (0 + 757) => x"00000000", (0 + 758) => x"00000000", (0 + 759) => x"00000000", (0 + 760) => x"00000000", (0 + 761) => x"00000000", (0 + 762) => x"00000000", (0 + 763) => x"00000000", (0 + 764) => x"00000000", (0 + 765) => x"00000000", (0 + 766) => x"00000000", (0 + 767) => x"00000000", (0 + 768) => x"00000000", (0 + 769) => x"00000000", (0 + 770) => x"00000000", (0 + 771) => x"00000000", (0 + 772) => x"00000000", (0 + 773) => x"00000000", (0 + 774) => x"00000000", (0 + 775) => x"00000000", (0 + 776) => x"00000000", (0 + 777) => x"00000000", (0 + 778) => x"00000000", (0 + 779) => x"00000000", (0 + 780) => x"00000000", (0 + 781) => x"00000000", (0 + 782) => x"00000000", (0 + 783) => x"00000000", (0 + 784) => x"00000000", (0 + 785) => x"00000000", (0 + 786) => x"00000000", (0 + 787) => x"00000000", (0 + 788) => x"00000000", (0 + 789) => x"00000000", (0 + 790) => x"00000000", (0 + 791) => x"00000000", (0 + 792) => x"00000000", (0 + 793) => x"00000000", (0 + 794) => x"00000000", (0 + 795) => x"00000000", (0 + 796) => x"00000000", (0 + 797) => x"00000000", (0 + 798) => x"00000000", (0 + 799) => x"00000000", (0 + 800) => x"00000000", (0 + 801) => x"00000000", (0 + 802) => x"00000000", (0 + 803) => x"00000000", (0 + 804) => x"00000000", (0 + 805) => x"00000000", (0 + 806) => x"00000000", (0 + 807) => x"00000000", (0 + 808) => x"00000000", (0 + 809) => x"00000000", (0 + 810) => x"00000000", (0 + 811) => x"00000000", (0 + 812) => x"00000000", (0 + 813) => x"00000000", (0 + 814) => x"00000000", (0 + 815) => x"00000000", (0 + 816) => x"00000000", (0 + 817) => x"00000000", (0 + 818) => x"00000000", (0 + 819) => x"00000000", (0 + 820) => x"00000000", (0 + 821) => x"00000000", (0 + 822) => x"00000000", (0 + 823) => x"00000000", (0 + 824) => x"00000000", (0 + 825) => x"00000000", (0 + 826) => x"00000000", (0 + 827) => x"00000000", (0 + 828) => x"00000000", (0 + 829) => x"00000000", (0 + 830) => x"00000000", (0 + 831) => x"00000000", (0 + 832) => x"00000000", (0 + 833) => x"00000000", (0 + 834) => x"00000000", (0 + 835) => x"00000000", (0 + 836) => x"00000000", (0 + 837) => x"00000000", (0 + 838) => x"00000000", (0 + 839) => x"00000000", (0 + 840) => x"00000000", (0 + 841) => x"00000000", (0 + 842) => x"00000000", (0 + 843) => x"00000000", (0 + 844) => x"00000000", (0 + 845) => x"00000000", (0 + 846) => x"00000000", (0 + 847) => x"00000000", (0 + 848) => x"00000000", (0 + 849) => x"00000000", (0 + 850) => x"00000000", (0 + 851) => x"00000000", (0 + 852) => x"00000000", (0 + 853) => x"00000000", (0 + 854) => x"00000000", (0 + 855) => x"00000000", (0 + 856) => x"00000000", (0 + 857) => x"00000000", (0 + 858) => x"00000000", (0 + 859) => x"00000000", (0 + 860) => x"00000000", (0 + 861) => x"00000000", (0 + 862) => x"00000000", (0 + 863) => x"00000000", (0 + 864) => x"00000000", (0 + 865) => x"00000000", (0 + 866) => x"00000000", (0 + 867) => x"00000000", (0 + 868) => x"00000000", (0 + 869) => x"00000000", (0 + 870) => x"00000000", (0 + 871) => x"00000000", (0 + 872) => x"00000000", (0 + 873) => x"00000000", (0 + 874) => x"00000000", (0 + 875) => x"00000000", (0 + 876) => x"00000000", (0 + 877) => x"00000000", (0 + 878) => x"00000000", (0 + 879) => x"00000000", (0 + 880) => x"00000000", (0 + 881) => x"00000000", (0 + 882) => x"00000000", (0 + 883) => x"00000000", (0 + 884) => x"00000000", (0 + 885) => x"00000000", (0 + 886) => x"00000000", (0 + 887) => x"00000000", (0 + 888) => x"00000000", (0 + 889) => x"00000000", (0 + 890) => x"00000000", (0 + 891) => x"00000000", (0 + 892) => x"00000000", (0 + 893) => x"00000000", (0 + 894) => x"00000000", (0 + 895) => x"00000000", (0 + 896) => x"00000000", (0 + 897) => x"00000000", (0 + 898) => x"00000000", (0 + 899) => x"00000000", (0 + 900) => x"00000000", (0 + 901) => x"00000000", (0 + 902) => x"00000000", (0 + 903) => x"00000000", (0 + 904) => x"00000000", (0 + 905) => x"00000000", (0 + 906) => x"00000000", (0 + 907) => x"00000000", (0 + 908) => x"00000000", (0 + 909) => x"00000000", (0 + 910) => x"00000000", (0 + 911) => x"00000000", (0 + 912) => x"00000000", (0 + 913) => x"00000000", (0 + 914) => x"00000000", (0 + 915) => x"00000000", (0 + 916) => x"00000000", (0 + 917) => x"00000000", (0 + 918) => x"00000000", (0 + 919) => x"00000000", (0 + 920) => x"00000000", (0 + 921) => x"00000000", (0 + 922) => x"00000000", (0 + 923) => x"00000000", (0 + 924) => x"00000000", (0 + 925) => x"00000000", (0 + 926) => x"00000000", (0 + 927) => x"00000000", (0 + 928) => x"00000000", (0 + 929) => x"00000000", (0 + 930) => x"00000000", (0 + 931) => x"00000000", (0 + 932) => x"00000000", (0 + 933) => x"00000000", (0 + 934) => x"00000000", (0 + 935) => x"00000000", (0 + 936) => x"00000000", (0 + 937) => x"00000000", (0 + 938) => x"00000000", (0 + 939) => x"00000000", (0 + 940) => x"00000000", (0 + 941) => x"00000000", (0 + 942) => x"00000000", (0 + 943) => x"00000000", (0 + 944) => x"00000000", (0 + 945) => x"00000000", (0 + 946) => x"00000000", (0 + 947) => x"00000000", (0 + 948) => x"00000000", (0 + 949) => x"00000000", (0 + 950) => x"00000000", (0 + 951) => x"00000000", (0 + 952) => x"00000000", (0 + 953) => x"00000000", (0 + 954) => x"00000000", (0 + 955) => x"00000000", (0 + 956) => x"00000000", (0 + 957) => x"00000000", (0 + 958) => x"00000000", (0 + 959) => x"00000000", (0 + 960) => x"00000000", (0 + 961) => x"00000000", (0 + 962) => x"00000000", (0 + 963) => x"00000000", (0 + 964) => x"00000000", (0 + 965) => x"00000000", (0 + 966) => x"00000000", (0 + 967) => x"00000000", (0 + 968) => x"00000000", (0 + 969) => x"00000000", (0 + 970) => x"00000000", (0 + 971) => x"00000000", (0 + 972) => x"00000000", (0 + 973) => x"00000000", (0 + 974) => x"00000000", (0 + 975) => x"00000000", (0 + 976) => x"00000000", (0 + 977) => x"00000000", (0 + 978) => x"00000000", (0 + 979) => x"00000000", (0 + 980) => x"00000000", (0 + 981) => x"00000000", (0 + 982) => x"00000000", (0 + 983) => x"00000000", (0 + 984) => x"00000000", (0 + 985) => x"00000000", (0 + 986) => x"00000000", (0 + 987) => x"00000000", (0 + 988) => x"00000000", (0 + 989) => x"00000000", (0 + 990) => x"00000000", (0 + 991) => x"00000000", (0 + 992) => x"00000000", (0 + 993) => x"00000000", (0 + 994) => x"00000000", (0 + 995) => x"00000000", (0 + 996) => x"00000000", (0 + 997) => x"00000000", (0 + 998) => x"00000000", (0 + 999) => x"00000000", (0 + 1000) => x"00000000", (0 + 1001) => x"00000000", (0 + 1002) => x"00000000", (0 + 1003) => x"00000000", (0 + 1004) => x"00000000", (0 + 1005) => x"00000000", (0 + 1006) => x"00000000", (0 + 1007) => x"00000000", (0 + 1008) => x"00000000", (0 + 1009) => x"00000000", (0 + 1010) => x"00000000", (0 + 1011) => x"00000000", (0 + 1012) => x"00000000", (0 + 1013) => x"00000000", (0 + 1014) => x"00000000", (0 + 1015) => x"00000000", (0 + 1016) => x"00000000", (0 + 1017) => x"00000000", (0 + 1018) => x"00000000", (0 + 1019) => x"00000000", (0 + 1020) => x"00000000", (0 + 1021) => x"00000000", (0 + 1022) => x"00000000", (0 + 1023) => x"00000000", 