(0 + 0) => x"17", (0 + 1) => x"01", (0 + 2) => x"00", (0 + 3) => x"00", (0 + 4) => x"13", (0 + 5) => x"01", (0 + 6) => x"01", (0 + 7) => x"0b", (0 + 8) => x"6f", (0 + 9) => x"00", (0 + 10) => x"40", (0 + 11) => x"00", (0 + 12) => x"13", (0 + 13) => x"01", (0 + 14) => x"01", (0 + 15) => x"ff", (0 + 16) => x"23", (0 + 17) => x"34", (0 + 18) => x"81", (0 + 19) => x"00", (0 + 20) => x"13", (0 + 21) => x"04", (0 + 22) => x"01", (0 + 23) => x"01", (0 + 24) => x"93", (0 + 25) => x"07", (0 + 26) => x"90", (0 + 27) => x"00", (0 + 28) => x"93", (0 + 29) => x"97", (0 + 30) => x"c7", (0 + 31) => x"01", (0 + 32) => x"13", (0 + 33) => x"07", (0 + 34) => x"f0", (0 + 35) => x"ff", (0 + 36) => x"23", (0 + 37) => x"90", (0 + 38) => x"e7", (0 + 39) => x"00", (0 + 40) => x"6f", (0 + 41) => x"00", (0 + 42) => x"00", (0 + 43) => x"00", (0 + 44) => x"00", 